module numbers_rom
	(
		input wire clk,
		input wire [7:0] row,
		input wire [3:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [7:0] row_reg;
	reg [3:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		12'b000000000000: color_data = 12'b111111111111;
		12'b000000000001: color_data = 12'b111111111111;
		12'b000000000010: color_data = 12'b111111111111;
		12'b000000000011: color_data = 12'b111111111111;
		12'b000000000100: color_data = 12'b111111111111;
		12'b000000000101: color_data = 12'b111111111111;
		12'b000000000110: color_data = 12'b111111111111;
		12'b000000000111: color_data = 12'b111111111111;
		12'b000000001000: color_data = 12'b111111111111;
		12'b000000001001: color_data = 12'b111111111111;
		12'b000000001010: color_data = 12'b111111111111;
		12'b000000001011: color_data = 12'b111111111111;
		12'b000000001100: color_data = 12'b111111111111;
		12'b000000001101: color_data = 12'b111111111111;
		12'b000000001110: color_data = 12'b111111111111;
		12'b000000001111: color_data = 12'b111111111111;

		12'b000000010000: color_data = 12'b111111111111;
		12'b000000010001: color_data = 12'b111111111111;
		12'b000000010010: color_data = 12'b111111111111;
		12'b000000010011: color_data = 12'b111111111111;
		12'b000000010100: color_data = 12'b000000000000;
		12'b000000010101: color_data = 12'b000000000000;
		12'b000000010110: color_data = 12'b000000000000;
		12'b000000010111: color_data = 12'b000000000000;
		12'b000000011000: color_data = 12'b000000000000;
		12'b000000011001: color_data = 12'b000000000000;
		12'b000000011010: color_data = 12'b000000000000;
		12'b000000011011: color_data = 12'b111111111111;
		12'b000000011100: color_data = 12'b111111111111;
		12'b000000011101: color_data = 12'b111111111111;
		12'b000000011110: color_data = 12'b111111111111;
		12'b000000011111: color_data = 12'b111111111111;

		12'b000000100000: color_data = 12'b111111111111;
		12'b000000100001: color_data = 12'b111111111111;
		12'b000000100010: color_data = 12'b111111111111;
		12'b000000100011: color_data = 12'b111111111111;
		12'b000000100100: color_data = 12'b000000000000;
		12'b000000100101: color_data = 12'b111111111111;
		12'b000000100110: color_data = 12'b111111111111;
		12'b000000100111: color_data = 12'b111111111111;
		12'b000000101000: color_data = 12'b111111111111;
		12'b000000101001: color_data = 12'b111111111111;
		12'b000000101010: color_data = 12'b000000000000;
		12'b000000101011: color_data = 12'b111111111111;
		12'b000000101100: color_data = 12'b111111111111;
		12'b000000101101: color_data = 12'b111111111111;
		12'b000000101110: color_data = 12'b111111111111;
		12'b000000101111: color_data = 12'b111111111111;

		12'b000000110000: color_data = 12'b111111111111;
		12'b000000110001: color_data = 12'b111111111111;
		12'b000000110010: color_data = 12'b111111111111;
		12'b000000110011: color_data = 12'b111111111111;
		12'b000000110100: color_data = 12'b000000000000;
		12'b000000110101: color_data = 12'b111111111111;
		12'b000000110110: color_data = 12'b111111111111;
		12'b000000110111: color_data = 12'b111111111111;
		12'b000000111000: color_data = 12'b111111111111;
		12'b000000111001: color_data = 12'b111111111111;
		12'b000000111010: color_data = 12'b000000000000;
		12'b000000111011: color_data = 12'b111111111111;
		12'b000000111100: color_data = 12'b111111111111;
		12'b000000111101: color_data = 12'b111111111111;
		12'b000000111110: color_data = 12'b111111111111;
		12'b000000111111: color_data = 12'b111111111111;

		12'b000001000000: color_data = 12'b111111111111;
		12'b000001000001: color_data = 12'b111111111111;
		12'b000001000010: color_data = 12'b111111111111;
		12'b000001000011: color_data = 12'b111111111111;
		12'b000001000100: color_data = 12'b000000000000;
		12'b000001000101: color_data = 12'b111111111111;
		12'b000001000110: color_data = 12'b111111111111;
		12'b000001000111: color_data = 12'b111111111111;
		12'b000001001000: color_data = 12'b111111111111;
		12'b000001001001: color_data = 12'b111111111111;
		12'b000001001010: color_data = 12'b000000000000;
		12'b000001001011: color_data = 12'b111111111111;
		12'b000001001100: color_data = 12'b111111111111;
		12'b000001001101: color_data = 12'b111111111111;
		12'b000001001110: color_data = 12'b111111111111;
		12'b000001001111: color_data = 12'b111111111111;

		12'b000001010000: color_data = 12'b111111111111;
		12'b000001010001: color_data = 12'b111111111111;
		12'b000001010010: color_data = 12'b111111111111;
		12'b000001010011: color_data = 12'b111111111111;
		12'b000001010100: color_data = 12'b000000000000;
		12'b000001010101: color_data = 12'b111111111111;
		12'b000001010110: color_data = 12'b111111111111;
		12'b000001010111: color_data = 12'b111111111111;
		12'b000001011000: color_data = 12'b111111111111;
		12'b000001011001: color_data = 12'b111111111111;
		12'b000001011010: color_data = 12'b000000000000;
		12'b000001011011: color_data = 12'b111111111111;
		12'b000001011100: color_data = 12'b111111111111;
		12'b000001011101: color_data = 12'b111111111111;
		12'b000001011110: color_data = 12'b111111111111;
		12'b000001011111: color_data = 12'b111111111111;

		12'b000001100000: color_data = 12'b111111111111;
		12'b000001100001: color_data = 12'b111111111111;
		12'b000001100010: color_data = 12'b111111111111;
		12'b000001100011: color_data = 12'b111111111111;
		12'b000001100100: color_data = 12'b000000000000;
		12'b000001100101: color_data = 12'b111111111111;
		12'b000001100110: color_data = 12'b111111111111;
		12'b000001100111: color_data = 12'b111111111111;
		12'b000001101000: color_data = 12'b111111111111;
		12'b000001101001: color_data = 12'b111111111111;
		12'b000001101010: color_data = 12'b000000000000;
		12'b000001101011: color_data = 12'b111111111111;
		12'b000001101100: color_data = 12'b111111111111;
		12'b000001101101: color_data = 12'b111111111111;
		12'b000001101110: color_data = 12'b111111111111;
		12'b000001101111: color_data = 12'b111111111111;

		12'b000001110000: color_data = 12'b111111111111;
		12'b000001110001: color_data = 12'b111111111111;
		12'b000001110010: color_data = 12'b111111111111;
		12'b000001110011: color_data = 12'b111111111111;
		12'b000001110100: color_data = 12'b000000000000;
		12'b000001110101: color_data = 12'b111111111111;
		12'b000001110110: color_data = 12'b111111111111;
		12'b000001110111: color_data = 12'b111111111111;
		12'b000001111000: color_data = 12'b111111111111;
		12'b000001111001: color_data = 12'b111111111111;
		12'b000001111010: color_data = 12'b000000000000;
		12'b000001111011: color_data = 12'b111111111111;
		12'b000001111100: color_data = 12'b111111111111;
		12'b000001111101: color_data = 12'b111111111111;
		12'b000001111110: color_data = 12'b111111111111;
		12'b000001111111: color_data = 12'b111111111111;

		12'b000010000000: color_data = 12'b111111111111;
		12'b000010000001: color_data = 12'b111111111111;
		12'b000010000010: color_data = 12'b111111111111;
		12'b000010000011: color_data = 12'b111111111111;
		12'b000010000100: color_data = 12'b000000000000;
		12'b000010000101: color_data = 12'b111111111111;
		12'b000010000110: color_data = 12'b111111111111;
		12'b000010000111: color_data = 12'b111111111111;
		12'b000010001000: color_data = 12'b111111111111;
		12'b000010001001: color_data = 12'b111111111111;
		12'b000010001010: color_data = 12'b000000000000;
		12'b000010001011: color_data = 12'b111111111111;
		12'b000010001100: color_data = 12'b111111111111;
		12'b000010001101: color_data = 12'b111111111111;
		12'b000010001110: color_data = 12'b111111111111;
		12'b000010001111: color_data = 12'b111111111111;

		12'b000010010000: color_data = 12'b111111111111;
		12'b000010010001: color_data = 12'b111111111111;
		12'b000010010010: color_data = 12'b111111111111;
		12'b000010010011: color_data = 12'b111111111111;
		12'b000010010100: color_data = 12'b000000000000;
		12'b000010010101: color_data = 12'b111111111111;
		12'b000010010110: color_data = 12'b111111111111;
		12'b000010010111: color_data = 12'b111111111111;
		12'b000010011000: color_data = 12'b111111111111;
		12'b000010011001: color_data = 12'b111111111111;
		12'b000010011010: color_data = 12'b000000000000;
		12'b000010011011: color_data = 12'b111111111111;
		12'b000010011100: color_data = 12'b111111111111;
		12'b000010011101: color_data = 12'b111111111111;
		12'b000010011110: color_data = 12'b111111111111;
		12'b000010011111: color_data = 12'b111111111111;

		12'b000010100000: color_data = 12'b111111111111;
		12'b000010100001: color_data = 12'b111111111111;
		12'b000010100010: color_data = 12'b111111111111;
		12'b000010100011: color_data = 12'b111111111111;
		12'b000010100100: color_data = 12'b000000000000;
		12'b000010100101: color_data = 12'b111111111111;
		12'b000010100110: color_data = 12'b111111111111;
		12'b000010100111: color_data = 12'b111111111111;
		12'b000010101000: color_data = 12'b111111111111;
		12'b000010101001: color_data = 12'b111111111111;
		12'b000010101010: color_data = 12'b000000000000;
		12'b000010101011: color_data = 12'b111111111111;
		12'b000010101100: color_data = 12'b111111111111;
		12'b000010101101: color_data = 12'b111111111111;
		12'b000010101110: color_data = 12'b111111111111;
		12'b000010101111: color_data = 12'b111111111111;

		12'b000010110000: color_data = 12'b111111111111;
		12'b000010110001: color_data = 12'b111111111111;
		12'b000010110010: color_data = 12'b111111111111;
		12'b000010110011: color_data = 12'b111111111111;
		12'b000010110100: color_data = 12'b000000000000;
		12'b000010110101: color_data = 12'b111111111111;
		12'b000010110110: color_data = 12'b111111111111;
		12'b000010110111: color_data = 12'b111111111111;
		12'b000010111000: color_data = 12'b111111111111;
		12'b000010111001: color_data = 12'b111111111111;
		12'b000010111010: color_data = 12'b000000000000;
		12'b000010111011: color_data = 12'b111111111111;
		12'b000010111100: color_data = 12'b111111111111;
		12'b000010111101: color_data = 12'b111111111111;
		12'b000010111110: color_data = 12'b111111111111;
		12'b000010111111: color_data = 12'b111111111111;

		12'b000011000000: color_data = 12'b111111111111;
		12'b000011000001: color_data = 12'b111111111111;
		12'b000011000010: color_data = 12'b111111111111;
		12'b000011000011: color_data = 12'b111111111111;
		12'b000011000100: color_data = 12'b000000000000;
		12'b000011000101: color_data = 12'b111111111111;
		12'b000011000110: color_data = 12'b111111111111;
		12'b000011000111: color_data = 12'b111111111111;
		12'b000011001000: color_data = 12'b111111111111;
		12'b000011001001: color_data = 12'b111111111111;
		12'b000011001010: color_data = 12'b000000000000;
		12'b000011001011: color_data = 12'b111111111111;
		12'b000011001100: color_data = 12'b111111111111;
		12'b000011001101: color_data = 12'b111111111111;
		12'b000011001110: color_data = 12'b111111111111;
		12'b000011001111: color_data = 12'b111111111111;

		12'b000011010000: color_data = 12'b111111111111;
		12'b000011010001: color_data = 12'b111111111111;
		12'b000011010010: color_data = 12'b111111111111;
		12'b000011010011: color_data = 12'b111111111111;
		12'b000011010100: color_data = 12'b000000000000;
		12'b000011010101: color_data = 12'b000000000000;
		12'b000011010110: color_data = 12'b000000000000;
		12'b000011010111: color_data = 12'b000000000000;
		12'b000011011000: color_data = 12'b000000000000;
		12'b000011011001: color_data = 12'b000000000000;
		12'b000011011010: color_data = 12'b000000000000;
		12'b000011011011: color_data = 12'b111111111111;
		12'b000011011100: color_data = 12'b111111111111;
		12'b000011011101: color_data = 12'b111111111111;
		12'b000011011110: color_data = 12'b111111111111;
		12'b000011011111: color_data = 12'b111111111111;

		12'b000011100000: color_data = 12'b111111111111;
		12'b000011100001: color_data = 12'b111111111111;
		12'b000011100010: color_data = 12'b111111111111;
		12'b000011100011: color_data = 12'b111111111111;
		12'b000011100100: color_data = 12'b111111111111;
		12'b000011100101: color_data = 12'b111111111111;
		12'b000011100110: color_data = 12'b111111111111;
		12'b000011100111: color_data = 12'b111111111111;
		12'b000011101000: color_data = 12'b111111111111;
		12'b000011101001: color_data = 12'b111111111111;
		12'b000011101010: color_data = 12'b111111111111;
		12'b000011101011: color_data = 12'b111111111111;
		12'b000011101100: color_data = 12'b111111111111;
		12'b000011101101: color_data = 12'b111111111111;
		12'b000011101110: color_data = 12'b111111111111;
		12'b000011101111: color_data = 12'b111111111111;

		12'b000011110000: color_data = 12'b111111111111;
		12'b000011110001: color_data = 12'b111111111111;
		12'b000011110010: color_data = 12'b111111111111;
		12'b000011110011: color_data = 12'b111111111111;
		12'b000011110100: color_data = 12'b111111111111;
		12'b000011110101: color_data = 12'b111111111111;
		12'b000011110110: color_data = 12'b111111111111;
		12'b000011110111: color_data = 12'b111111111111;
		12'b000011111000: color_data = 12'b111111111111;
		12'b000011111001: color_data = 12'b111111111111;
		12'b000011111010: color_data = 12'b111111111111;
		12'b000011111011: color_data = 12'b111111111111;
		12'b000011111100: color_data = 12'b111111111111;
		12'b000011111101: color_data = 12'b111111111111;
		12'b000011111110: color_data = 12'b111111111111;
		12'b000011111111: color_data = 12'b111111111111;

		12'b000100000000: color_data = 12'b111111111111;
		12'b000100000001: color_data = 12'b111111111111;
		12'b000100000010: color_data = 12'b111111111111;
		12'b000100000011: color_data = 12'b111111111111;
		12'b000100000100: color_data = 12'b111111111111;
		12'b000100000101: color_data = 12'b111111111111;
		12'b000100000110: color_data = 12'b111111111111;
		12'b000100000111: color_data = 12'b111111111111;
		12'b000100001000: color_data = 12'b111111111111;
		12'b000100001001: color_data = 12'b111111111111;
		12'b000100001010: color_data = 12'b111111111111;
		12'b000100001011: color_data = 12'b111111111111;
		12'b000100001100: color_data = 12'b111111111111;
		12'b000100001101: color_data = 12'b111111111111;
		12'b000100001110: color_data = 12'b111111111111;
		12'b000100001111: color_data = 12'b111111111111;

		12'b000100010000: color_data = 12'b111111111111;
		12'b000100010001: color_data = 12'b111111111111;
		12'b000100010010: color_data = 12'b111111111111;
		12'b000100010011: color_data = 12'b111111111111;
		12'b000100010100: color_data = 12'b111111111111;
		12'b000100010101: color_data = 12'b111111111111;
		12'b000100010110: color_data = 12'b000000000000;
		12'b000100010111: color_data = 12'b000000000000;
		12'b000100011000: color_data = 12'b111111111111;
		12'b000100011001: color_data = 12'b111111111111;
		12'b000100011010: color_data = 12'b111111111111;
		12'b000100011011: color_data = 12'b111111111111;
		12'b000100011100: color_data = 12'b111111111111;
		12'b000100011101: color_data = 12'b111111111111;
		12'b000100011110: color_data = 12'b111111111111;
		12'b000100011111: color_data = 12'b111111111111;

		12'b000100100000: color_data = 12'b111111111111;
		12'b000100100001: color_data = 12'b111111111111;
		12'b000100100010: color_data = 12'b111111111111;
		12'b000100100011: color_data = 12'b111111111111;
		12'b000100100100: color_data = 12'b111111111111;
		12'b000100100101: color_data = 12'b000000000000;
		12'b000100100110: color_data = 12'b000000000000;
		12'b000100100111: color_data = 12'b000000000000;
		12'b000100101000: color_data = 12'b111111111111;
		12'b000100101001: color_data = 12'b111111111111;
		12'b000100101010: color_data = 12'b111111111111;
		12'b000100101011: color_data = 12'b111111111111;
		12'b000100101100: color_data = 12'b111111111111;
		12'b000100101101: color_data = 12'b111111111111;
		12'b000100101110: color_data = 12'b111111111111;
		12'b000100101111: color_data = 12'b111111111111;

		12'b000100110000: color_data = 12'b111111111111;
		12'b000100110001: color_data = 12'b111111111111;
		12'b000100110010: color_data = 12'b111111111111;
		12'b000100110011: color_data = 12'b111111111111;
		12'b000100110100: color_data = 12'b000000000000;
		12'b000100110101: color_data = 12'b000000000000;
		12'b000100110110: color_data = 12'b111111111111;
		12'b000100110111: color_data = 12'b000000000000;
		12'b000100111000: color_data = 12'b111111111111;
		12'b000100111001: color_data = 12'b111111111111;
		12'b000100111010: color_data = 12'b111111111111;
		12'b000100111011: color_data = 12'b111111111111;
		12'b000100111100: color_data = 12'b111111111111;
		12'b000100111101: color_data = 12'b111111111111;
		12'b000100111110: color_data = 12'b111111111111;
		12'b000100111111: color_data = 12'b111111111111;

		12'b000101000000: color_data = 12'b111111111111;
		12'b000101000001: color_data = 12'b111111111111;
		12'b000101000010: color_data = 12'b111111111111;
		12'b000101000011: color_data = 12'b111111111111;
		12'b000101000100: color_data = 12'b000000000000;
		12'b000101000101: color_data = 12'b111111111111;
		12'b000101000110: color_data = 12'b111111111111;
		12'b000101000111: color_data = 12'b000000000000;
		12'b000101001000: color_data = 12'b111111111111;
		12'b000101001001: color_data = 12'b111111111111;
		12'b000101001010: color_data = 12'b111111111111;
		12'b000101001011: color_data = 12'b111111111111;
		12'b000101001100: color_data = 12'b111111111111;
		12'b000101001101: color_data = 12'b111111111111;
		12'b000101001110: color_data = 12'b111111111111;
		12'b000101001111: color_data = 12'b111111111111;

		12'b000101010000: color_data = 12'b111111111111;
		12'b000101010001: color_data = 12'b111111111111;
		12'b000101010010: color_data = 12'b111111111111;
		12'b000101010011: color_data = 12'b111111111111;
		12'b000101010100: color_data = 12'b111111111111;
		12'b000101010101: color_data = 12'b111111111111;
		12'b000101010110: color_data = 12'b111111111111;
		12'b000101010111: color_data = 12'b000000000000;
		12'b000101011000: color_data = 12'b111111111111;
		12'b000101011001: color_data = 12'b111111111111;
		12'b000101011010: color_data = 12'b111111111111;
		12'b000101011011: color_data = 12'b111111111111;
		12'b000101011100: color_data = 12'b111111111111;
		12'b000101011101: color_data = 12'b111111111111;
		12'b000101011110: color_data = 12'b111111111111;
		12'b000101011111: color_data = 12'b111111111111;

		12'b000101100000: color_data = 12'b111111111111;
		12'b000101100001: color_data = 12'b111111111111;
		12'b000101100010: color_data = 12'b111111111111;
		12'b000101100011: color_data = 12'b111111111111;
		12'b000101100100: color_data = 12'b111111111111;
		12'b000101100101: color_data = 12'b111111111111;
		12'b000101100110: color_data = 12'b111111111111;
		12'b000101100111: color_data = 12'b000000000000;
		12'b000101101000: color_data = 12'b111111111111;
		12'b000101101001: color_data = 12'b111111111111;
		12'b000101101010: color_data = 12'b111111111111;
		12'b000101101011: color_data = 12'b111111111111;
		12'b000101101100: color_data = 12'b111111111111;
		12'b000101101101: color_data = 12'b111111111111;
		12'b000101101110: color_data = 12'b111111111111;
		12'b000101101111: color_data = 12'b111111111111;

		12'b000101110000: color_data = 12'b111111111111;
		12'b000101110001: color_data = 12'b111111111111;
		12'b000101110010: color_data = 12'b111111111111;
		12'b000101110011: color_data = 12'b111111111111;
		12'b000101110100: color_data = 12'b111111111111;
		12'b000101110101: color_data = 12'b111111111111;
		12'b000101110110: color_data = 12'b111111111111;
		12'b000101110111: color_data = 12'b000000000000;
		12'b000101111000: color_data = 12'b111111111111;
		12'b000101111001: color_data = 12'b111111111111;
		12'b000101111010: color_data = 12'b111111111111;
		12'b000101111011: color_data = 12'b111111111111;
		12'b000101111100: color_data = 12'b111111111111;
		12'b000101111101: color_data = 12'b111111111111;
		12'b000101111110: color_data = 12'b111111111111;
		12'b000101111111: color_data = 12'b111111111111;

		12'b000110000000: color_data = 12'b111111111111;
		12'b000110000001: color_data = 12'b111111111111;
		12'b000110000010: color_data = 12'b111111111111;
		12'b000110000011: color_data = 12'b111111111111;
		12'b000110000100: color_data = 12'b111111111111;
		12'b000110000101: color_data = 12'b111111111111;
		12'b000110000110: color_data = 12'b111111111111;
		12'b000110000111: color_data = 12'b000000000000;
		12'b000110001000: color_data = 12'b111111111111;
		12'b000110001001: color_data = 12'b111111111111;
		12'b000110001010: color_data = 12'b111111111111;
		12'b000110001011: color_data = 12'b111111111111;
		12'b000110001100: color_data = 12'b111111111111;
		12'b000110001101: color_data = 12'b111111111111;
		12'b000110001110: color_data = 12'b111111111111;
		12'b000110001111: color_data = 12'b111111111111;

		12'b000110010000: color_data = 12'b111111111111;
		12'b000110010001: color_data = 12'b111111111111;
		12'b000110010010: color_data = 12'b111111111111;
		12'b000110010011: color_data = 12'b111111111111;
		12'b000110010100: color_data = 12'b111111111111;
		12'b000110010101: color_data = 12'b111111111111;
		12'b000110010110: color_data = 12'b111111111111;
		12'b000110010111: color_data = 12'b000000000000;
		12'b000110011000: color_data = 12'b111111111111;
		12'b000110011001: color_data = 12'b111111111111;
		12'b000110011010: color_data = 12'b111111111111;
		12'b000110011011: color_data = 12'b111111111111;
		12'b000110011100: color_data = 12'b111111111111;
		12'b000110011101: color_data = 12'b111111111111;
		12'b000110011110: color_data = 12'b111111111111;
		12'b000110011111: color_data = 12'b111111111111;

		12'b000110100000: color_data = 12'b111111111111;
		12'b000110100001: color_data = 12'b111111111111;
		12'b000110100010: color_data = 12'b111111111111;
		12'b000110100011: color_data = 12'b111111111111;
		12'b000110100100: color_data = 12'b111111111111;
		12'b000110100101: color_data = 12'b111111111111;
		12'b000110100110: color_data = 12'b111111111111;
		12'b000110100111: color_data = 12'b000000000000;
		12'b000110101000: color_data = 12'b111111111111;
		12'b000110101001: color_data = 12'b111111111111;
		12'b000110101010: color_data = 12'b111111111111;
		12'b000110101011: color_data = 12'b111111111111;
		12'b000110101100: color_data = 12'b111111111111;
		12'b000110101101: color_data = 12'b111111111111;
		12'b000110101110: color_data = 12'b111111111111;
		12'b000110101111: color_data = 12'b111111111111;

		12'b000110110000: color_data = 12'b111111111111;
		12'b000110110001: color_data = 12'b111111111111;
		12'b000110110010: color_data = 12'b111111111111;
		12'b000110110011: color_data = 12'b111111111111;
		12'b000110110100: color_data = 12'b111111111111;
		12'b000110110101: color_data = 12'b111111111111;
		12'b000110110110: color_data = 12'b111111111111;
		12'b000110110111: color_data = 12'b000000000000;
		12'b000110111000: color_data = 12'b111111111111;
		12'b000110111001: color_data = 12'b111111111111;
		12'b000110111010: color_data = 12'b111111111111;
		12'b000110111011: color_data = 12'b111111111111;
		12'b000110111100: color_data = 12'b111111111111;
		12'b000110111101: color_data = 12'b111111111111;
		12'b000110111110: color_data = 12'b111111111111;
		12'b000110111111: color_data = 12'b111111111111;

		12'b000111000000: color_data = 12'b111111111111;
		12'b000111000001: color_data = 12'b111111111111;
		12'b000111000010: color_data = 12'b111111111111;
		12'b000111000011: color_data = 12'b111111111111;
		12'b000111000100: color_data = 12'b111111111111;
		12'b000111000101: color_data = 12'b111111111111;
		12'b000111000110: color_data = 12'b111111111111;
		12'b000111000111: color_data = 12'b000000000000;
		12'b000111001000: color_data = 12'b111111111111;
		12'b000111001001: color_data = 12'b111111111111;
		12'b000111001010: color_data = 12'b111111111111;
		12'b000111001011: color_data = 12'b111111111111;
		12'b000111001100: color_data = 12'b111111111111;
		12'b000111001101: color_data = 12'b111111111111;
		12'b000111001110: color_data = 12'b111111111111;
		12'b000111001111: color_data = 12'b111111111111;

		12'b000111010000: color_data = 12'b111111111111;
		12'b000111010001: color_data = 12'b111111111111;
		12'b000111010010: color_data = 12'b111111111111;
		12'b000111010011: color_data = 12'b111111111111;
		12'b000111010100: color_data = 12'b000000000000;
		12'b000111010101: color_data = 12'b000000000000;
		12'b000111010110: color_data = 12'b000000000000;
		12'b000111010111: color_data = 12'b000000000000;
		12'b000111011000: color_data = 12'b000000000000;
		12'b000111011001: color_data = 12'b000000000000;
		12'b000111011010: color_data = 12'b000000000000;
		12'b000111011011: color_data = 12'b111111111111;
		12'b000111011100: color_data = 12'b111111111111;
		12'b000111011101: color_data = 12'b111111111111;
		12'b000111011110: color_data = 12'b111111111111;
		12'b000111011111: color_data = 12'b111111111111;

		12'b000111100000: color_data = 12'b111111111111;
		12'b000111100001: color_data = 12'b111111111111;
		12'b000111100010: color_data = 12'b111111111111;
		12'b000111100011: color_data = 12'b111111111111;
		12'b000111100100: color_data = 12'b111111111111;
		12'b000111100101: color_data = 12'b111111111111;
		12'b000111100110: color_data = 12'b111111111111;
		12'b000111100111: color_data = 12'b111111111111;
		12'b000111101000: color_data = 12'b111111111111;
		12'b000111101001: color_data = 12'b111111111111;
		12'b000111101010: color_data = 12'b111111111111;
		12'b000111101011: color_data = 12'b111111111111;
		12'b000111101100: color_data = 12'b111111111111;
		12'b000111101101: color_data = 12'b111111111111;
		12'b000111101110: color_data = 12'b111111111111;
		12'b000111101111: color_data = 12'b111111111111;

		12'b000111110000: color_data = 12'b111111111111;
		12'b000111110001: color_data = 12'b111111111111;
		12'b000111110010: color_data = 12'b111111111111;
		12'b000111110011: color_data = 12'b111111111111;
		12'b000111110100: color_data = 12'b111111111111;
		12'b000111110101: color_data = 12'b111111111111;
		12'b000111110110: color_data = 12'b111111111111;
		12'b000111110111: color_data = 12'b111111111111;
		12'b000111111000: color_data = 12'b111111111111;
		12'b000111111001: color_data = 12'b111111111111;
		12'b000111111010: color_data = 12'b111111111111;
		12'b000111111011: color_data = 12'b111111111111;
		12'b000111111100: color_data = 12'b111111111111;
		12'b000111111101: color_data = 12'b111111111111;
		12'b000111111110: color_data = 12'b111111111111;
		12'b000111111111: color_data = 12'b111111111111;

		12'b001000000000: color_data = 12'b111111111111;
		12'b001000000001: color_data = 12'b111111111111;
		12'b001000000010: color_data = 12'b111111111111;
		12'b001000000011: color_data = 12'b111111111111;
		12'b001000000100: color_data = 12'b111111111111;
		12'b001000000101: color_data = 12'b111111111111;
		12'b001000000110: color_data = 12'b111111111111;
		12'b001000000111: color_data = 12'b111111111111;
		12'b001000001000: color_data = 12'b111111111111;
		12'b001000001001: color_data = 12'b111111111111;
		12'b001000001010: color_data = 12'b111111111111;
		12'b001000001011: color_data = 12'b111111111111;
		12'b001000001100: color_data = 12'b111111111111;
		12'b001000001101: color_data = 12'b111111111111;
		12'b001000001110: color_data = 12'b111111111111;
		12'b001000001111: color_data = 12'b111111111111;

		12'b001000010000: color_data = 12'b111111111111;
		12'b001000010001: color_data = 12'b111111111111;
		12'b001000010010: color_data = 12'b111111111111;
		12'b001000010011: color_data = 12'b111111111111;
		12'b001000010100: color_data = 12'b000000000000;
		12'b001000010101: color_data = 12'b000000000000;
		12'b001000010110: color_data = 12'b000000000000;
		12'b001000010111: color_data = 12'b000000000000;
		12'b001000011000: color_data = 12'b000000000000;
		12'b001000011001: color_data = 12'b000000000000;
		12'b001000011010: color_data = 12'b000000000000;
		12'b001000011011: color_data = 12'b111111111111;
		12'b001000011100: color_data = 12'b111111111111;
		12'b001000011101: color_data = 12'b111111111111;
		12'b001000011110: color_data = 12'b111111111111;
		12'b001000011111: color_data = 12'b111111111111;

		12'b001000100000: color_data = 12'b111111111111;
		12'b001000100001: color_data = 12'b111111111111;
		12'b001000100010: color_data = 12'b111111111111;
		12'b001000100011: color_data = 12'b111111111111;
		12'b001000100100: color_data = 12'b000000000000;
		12'b001000100101: color_data = 12'b111111111111;
		12'b001000100110: color_data = 12'b111111111111;
		12'b001000100111: color_data = 12'b111111111111;
		12'b001000101000: color_data = 12'b111111111111;
		12'b001000101001: color_data = 12'b111111111111;
		12'b001000101010: color_data = 12'b000000000000;
		12'b001000101011: color_data = 12'b111111111111;
		12'b001000101100: color_data = 12'b111111111111;
		12'b001000101101: color_data = 12'b111111111111;
		12'b001000101110: color_data = 12'b111111111111;
		12'b001000101111: color_data = 12'b111111111111;

		12'b001000110000: color_data = 12'b111111111111;
		12'b001000110001: color_data = 12'b111111111111;
		12'b001000110010: color_data = 12'b111111111111;
		12'b001000110011: color_data = 12'b111111111111;
		12'b001000110100: color_data = 12'b000000000000;
		12'b001000110101: color_data = 12'b111111111111;
		12'b001000110110: color_data = 12'b111111111111;
		12'b001000110111: color_data = 12'b111111111111;
		12'b001000111000: color_data = 12'b111111111111;
		12'b001000111001: color_data = 12'b111111111111;
		12'b001000111010: color_data = 12'b000000000000;
		12'b001000111011: color_data = 12'b111111111111;
		12'b001000111100: color_data = 12'b111111111111;
		12'b001000111101: color_data = 12'b111111111111;
		12'b001000111110: color_data = 12'b111111111111;
		12'b001000111111: color_data = 12'b111111111111;

		12'b001001000000: color_data = 12'b111111111111;
		12'b001001000001: color_data = 12'b111111111111;
		12'b001001000010: color_data = 12'b111111111111;
		12'b001001000011: color_data = 12'b111111111111;
		12'b001001000100: color_data = 12'b000000000000;
		12'b001001000101: color_data = 12'b111111111111;
		12'b001001000110: color_data = 12'b111111111111;
		12'b001001000111: color_data = 12'b111111111111;
		12'b001001001000: color_data = 12'b111111111111;
		12'b001001001001: color_data = 12'b111111111111;
		12'b001001001010: color_data = 12'b000000000000;
		12'b001001001011: color_data = 12'b111111111111;
		12'b001001001100: color_data = 12'b111111111111;
		12'b001001001101: color_data = 12'b111111111111;
		12'b001001001110: color_data = 12'b111111111111;
		12'b001001001111: color_data = 12'b111111111111;

		12'b001001010000: color_data = 12'b111111111111;
		12'b001001010001: color_data = 12'b111111111111;
		12'b001001010010: color_data = 12'b111111111111;
		12'b001001010011: color_data = 12'b111111111111;
		12'b001001010100: color_data = 12'b000000000000;
		12'b001001010101: color_data = 12'b111111111111;
		12'b001001010110: color_data = 12'b111111111111;
		12'b001001010111: color_data = 12'b111111111111;
		12'b001001011000: color_data = 12'b111111111111;
		12'b001001011001: color_data = 12'b111111111111;
		12'b001001011010: color_data = 12'b000000000000;
		12'b001001011011: color_data = 12'b111111111111;
		12'b001001011100: color_data = 12'b111111111111;
		12'b001001011101: color_data = 12'b111111111111;
		12'b001001011110: color_data = 12'b111111111111;
		12'b001001011111: color_data = 12'b111111111111;

		12'b001001100000: color_data = 12'b111111111111;
		12'b001001100001: color_data = 12'b111111111111;
		12'b001001100010: color_data = 12'b111111111111;
		12'b001001100011: color_data = 12'b111111111111;
		12'b001001100100: color_data = 12'b111111111111;
		12'b001001100101: color_data = 12'b111111111111;
		12'b001001100110: color_data = 12'b111111111111;
		12'b001001100111: color_data = 12'b111111111111;
		12'b001001101000: color_data = 12'b111111111111;
		12'b001001101001: color_data = 12'b111111111111;
		12'b001001101010: color_data = 12'b000000000000;
		12'b001001101011: color_data = 12'b111111111111;
		12'b001001101100: color_data = 12'b111111111111;
		12'b001001101101: color_data = 12'b111111111111;
		12'b001001101110: color_data = 12'b111111111111;
		12'b001001101111: color_data = 12'b111111111111;

		12'b001001110000: color_data = 12'b111111111111;
		12'b001001110001: color_data = 12'b111111111111;
		12'b001001110010: color_data = 12'b111111111111;
		12'b001001110011: color_data = 12'b111111111111;
		12'b001001110100: color_data = 12'b111111111111;
		12'b001001110101: color_data = 12'b111111111111;
		12'b001001110110: color_data = 12'b111111111111;
		12'b001001110111: color_data = 12'b111111111111;
		12'b001001111000: color_data = 12'b111111111111;
		12'b001001111001: color_data = 12'b111111111111;
		12'b001001111010: color_data = 12'b000000000000;
		12'b001001111011: color_data = 12'b111111111111;
		12'b001001111100: color_data = 12'b111111111111;
		12'b001001111101: color_data = 12'b111111111111;
		12'b001001111110: color_data = 12'b111111111111;
		12'b001001111111: color_data = 12'b111111111111;

		12'b001010000000: color_data = 12'b111111111111;
		12'b001010000001: color_data = 12'b111111111111;
		12'b001010000010: color_data = 12'b111111111111;
		12'b001010000011: color_data = 12'b111111111111;
		12'b001010000100: color_data = 12'b111111111111;
		12'b001010000101: color_data = 12'b111111111111;
		12'b001010000110: color_data = 12'b111111111111;
		12'b001010000111: color_data = 12'b111111111111;
		12'b001010001000: color_data = 12'b111111111111;
		12'b001010001001: color_data = 12'b111111111111;
		12'b001010001010: color_data = 12'b000000000000;
		12'b001010001011: color_data = 12'b111111111111;
		12'b001010001100: color_data = 12'b111111111111;
		12'b001010001101: color_data = 12'b111111111111;
		12'b001010001110: color_data = 12'b111111111111;
		12'b001010001111: color_data = 12'b111111111111;

		12'b001010010000: color_data = 12'b111111111111;
		12'b001010010001: color_data = 12'b111111111111;
		12'b001010010010: color_data = 12'b111111111111;
		12'b001010010011: color_data = 12'b111111111111;
		12'b001010010100: color_data = 12'b000000000000;
		12'b001010010101: color_data = 12'b000000000000;
		12'b001010010110: color_data = 12'b000000000000;
		12'b001010010111: color_data = 12'b000000000000;
		12'b001010011000: color_data = 12'b000000000000;
		12'b001010011001: color_data = 12'b000000000000;
		12'b001010011010: color_data = 12'b000000000000;
		12'b001010011011: color_data = 12'b111111111111;
		12'b001010011100: color_data = 12'b111111111111;
		12'b001010011101: color_data = 12'b111111111111;
		12'b001010011110: color_data = 12'b111111111111;
		12'b001010011111: color_data = 12'b111111111111;

		12'b001010100000: color_data = 12'b111111111111;
		12'b001010100001: color_data = 12'b111111111111;
		12'b001010100010: color_data = 12'b111111111111;
		12'b001010100011: color_data = 12'b111111111111;
		12'b001010100100: color_data = 12'b000000000000;
		12'b001010100101: color_data = 12'b111111111111;
		12'b001010100110: color_data = 12'b111111111111;
		12'b001010100111: color_data = 12'b111111111111;
		12'b001010101000: color_data = 12'b111111111111;
		12'b001010101001: color_data = 12'b111111111111;
		12'b001010101010: color_data = 12'b111111111111;
		12'b001010101011: color_data = 12'b111111111111;
		12'b001010101100: color_data = 12'b111111111111;
		12'b001010101101: color_data = 12'b111111111111;
		12'b001010101110: color_data = 12'b111111111111;
		12'b001010101111: color_data = 12'b111111111111;

		12'b001010110000: color_data = 12'b111111111111;
		12'b001010110001: color_data = 12'b111111111111;
		12'b001010110010: color_data = 12'b111111111111;
		12'b001010110011: color_data = 12'b111111111111;
		12'b001010110100: color_data = 12'b000000000000;
		12'b001010110101: color_data = 12'b111111111111;
		12'b001010110110: color_data = 12'b111111111111;
		12'b001010110111: color_data = 12'b111111111111;
		12'b001010111000: color_data = 12'b111111111111;
		12'b001010111001: color_data = 12'b111111111111;
		12'b001010111010: color_data = 12'b111111111111;
		12'b001010111011: color_data = 12'b111111111111;
		12'b001010111100: color_data = 12'b111111111111;
		12'b001010111101: color_data = 12'b111111111111;
		12'b001010111110: color_data = 12'b111111111111;
		12'b001010111111: color_data = 12'b111111111111;

		12'b001011000000: color_data = 12'b111111111111;
		12'b001011000001: color_data = 12'b111111111111;
		12'b001011000010: color_data = 12'b111111111111;
		12'b001011000011: color_data = 12'b111111111111;
		12'b001011000100: color_data = 12'b000000000000;
		12'b001011000101: color_data = 12'b111111111111;
		12'b001011000110: color_data = 12'b111111111111;
		12'b001011000111: color_data = 12'b111111111111;
		12'b001011001000: color_data = 12'b111111111111;
		12'b001011001001: color_data = 12'b111111111111;
		12'b001011001010: color_data = 12'b111111111111;
		12'b001011001011: color_data = 12'b111111111111;
		12'b001011001100: color_data = 12'b111111111111;
		12'b001011001101: color_data = 12'b111111111111;
		12'b001011001110: color_data = 12'b111111111111;
		12'b001011001111: color_data = 12'b111111111111;

		12'b001011010000: color_data = 12'b111111111111;
		12'b001011010001: color_data = 12'b111111111111;
		12'b001011010010: color_data = 12'b111111111111;
		12'b001011010011: color_data = 12'b111111111111;
		12'b001011010100: color_data = 12'b000000000000;
		12'b001011010101: color_data = 12'b000000000000;
		12'b001011010110: color_data = 12'b000000000000;
		12'b001011010111: color_data = 12'b000000000000;
		12'b001011011000: color_data = 12'b000000000000;
		12'b001011011001: color_data = 12'b000000000000;
		12'b001011011010: color_data = 12'b000000000000;
		12'b001011011011: color_data = 12'b111111111111;
		12'b001011011100: color_data = 12'b111111111111;
		12'b001011011101: color_data = 12'b111111111111;
		12'b001011011110: color_data = 12'b111111111111;
		12'b001011011111: color_data = 12'b111111111111;

		12'b001011100000: color_data = 12'b111111111111;
		12'b001011100001: color_data = 12'b111111111111;
		12'b001011100010: color_data = 12'b111111111111;
		12'b001011100011: color_data = 12'b111111111111;
		12'b001011100100: color_data = 12'b111111111111;
		12'b001011100101: color_data = 12'b111111111111;
		12'b001011100110: color_data = 12'b111111111111;
		12'b001011100111: color_data = 12'b111111111111;
		12'b001011101000: color_data = 12'b111111111111;
		12'b001011101001: color_data = 12'b111111111111;
		12'b001011101010: color_data = 12'b111111111111;
		12'b001011101011: color_data = 12'b111111111111;
		12'b001011101100: color_data = 12'b111111111111;
		12'b001011101101: color_data = 12'b111111111111;
		12'b001011101110: color_data = 12'b111111111111;
		12'b001011101111: color_data = 12'b111111111111;

		12'b001011110000: color_data = 12'b111111111111;
		12'b001011110001: color_data = 12'b111111111111;
		12'b001011110010: color_data = 12'b111111111111;
		12'b001011110011: color_data = 12'b111111111111;
		12'b001011110100: color_data = 12'b111111111111;
		12'b001011110101: color_data = 12'b111111111111;
		12'b001011110110: color_data = 12'b111111111111;
		12'b001011110111: color_data = 12'b111111111111;
		12'b001011111000: color_data = 12'b111111111111;
		12'b001011111001: color_data = 12'b111111111111;
		12'b001011111010: color_data = 12'b111111111111;
		12'b001011111011: color_data = 12'b111111111111;
		12'b001011111100: color_data = 12'b111111111111;
		12'b001011111101: color_data = 12'b111111111111;
		12'b001011111110: color_data = 12'b111111111111;
		12'b001011111111: color_data = 12'b111111111111;

		12'b001100000000: color_data = 12'b111111111111;
		12'b001100000001: color_data = 12'b111111111111;
		12'b001100000010: color_data = 12'b111111111111;
		12'b001100000011: color_data = 12'b111111111111;
		12'b001100000100: color_data = 12'b111111111111;
		12'b001100000101: color_data = 12'b111111111111;
		12'b001100000110: color_data = 12'b111111111111;
		12'b001100000111: color_data = 12'b111111111111;
		12'b001100001000: color_data = 12'b111111111111;
		12'b001100001001: color_data = 12'b111111111111;
		12'b001100001010: color_data = 12'b111111111111;
		12'b001100001011: color_data = 12'b111111111111;
		12'b001100001100: color_data = 12'b111111111111;
		12'b001100001101: color_data = 12'b111111111111;
		12'b001100001110: color_data = 12'b111111111111;
		12'b001100001111: color_data = 12'b111111111111;

		12'b001100010000: color_data = 12'b111111111111;
		12'b001100010001: color_data = 12'b111111111111;
		12'b001100010010: color_data = 12'b111111111111;
		12'b001100010011: color_data = 12'b111111111111;
		12'b001100010100: color_data = 12'b000000000000;
		12'b001100010101: color_data = 12'b000000000000;
		12'b001100010110: color_data = 12'b000000000000;
		12'b001100010111: color_data = 12'b000000000000;
		12'b001100011000: color_data = 12'b000000000000;
		12'b001100011001: color_data = 12'b000000000000;
		12'b001100011010: color_data = 12'b000000000000;
		12'b001100011011: color_data = 12'b111111111111;
		12'b001100011100: color_data = 12'b111111111111;
		12'b001100011101: color_data = 12'b111111111111;
		12'b001100011110: color_data = 12'b111111111111;
		12'b001100011111: color_data = 12'b111111111111;

		12'b001100100000: color_data = 12'b111111111111;
		12'b001100100001: color_data = 12'b111111111111;
		12'b001100100010: color_data = 12'b111111111111;
		12'b001100100011: color_data = 12'b111111111111;
		12'b001100100100: color_data = 12'b000000000000;
		12'b001100100101: color_data = 12'b111111111111;
		12'b001100100110: color_data = 12'b111111111111;
		12'b001100100111: color_data = 12'b111111111111;
		12'b001100101000: color_data = 12'b111111111111;
		12'b001100101001: color_data = 12'b111111111111;
		12'b001100101010: color_data = 12'b000000000000;
		12'b001100101011: color_data = 12'b111111111111;
		12'b001100101100: color_data = 12'b111111111111;
		12'b001100101101: color_data = 12'b111111111111;
		12'b001100101110: color_data = 12'b111111111111;
		12'b001100101111: color_data = 12'b111111111111;

		12'b001100110000: color_data = 12'b111111111111;
		12'b001100110001: color_data = 12'b111111111111;
		12'b001100110010: color_data = 12'b111111111111;
		12'b001100110011: color_data = 12'b111111111111;
		12'b001100110100: color_data = 12'b000000000000;
		12'b001100110101: color_data = 12'b111111111111;
		12'b001100110110: color_data = 12'b111111111111;
		12'b001100110111: color_data = 12'b111111111111;
		12'b001100111000: color_data = 12'b111111111111;
		12'b001100111001: color_data = 12'b111111111111;
		12'b001100111010: color_data = 12'b000000000000;
		12'b001100111011: color_data = 12'b111111111111;
		12'b001100111100: color_data = 12'b111111111111;
		12'b001100111101: color_data = 12'b111111111111;
		12'b001100111110: color_data = 12'b111111111111;
		12'b001100111111: color_data = 12'b111111111111;

		12'b001101000000: color_data = 12'b111111111111;
		12'b001101000001: color_data = 12'b111111111111;
		12'b001101000010: color_data = 12'b111111111111;
		12'b001101000011: color_data = 12'b111111111111;
		12'b001101000100: color_data = 12'b000000000000;
		12'b001101000101: color_data = 12'b111111111111;
		12'b001101000110: color_data = 12'b111111111111;
		12'b001101000111: color_data = 12'b111111111111;
		12'b001101001000: color_data = 12'b111111111111;
		12'b001101001001: color_data = 12'b111111111111;
		12'b001101001010: color_data = 12'b000000000000;
		12'b001101001011: color_data = 12'b111111111111;
		12'b001101001100: color_data = 12'b111111111111;
		12'b001101001101: color_data = 12'b111111111111;
		12'b001101001110: color_data = 12'b111111111111;
		12'b001101001111: color_data = 12'b111111111111;

		12'b001101010000: color_data = 12'b111111111111;
		12'b001101010001: color_data = 12'b111111111111;
		12'b001101010010: color_data = 12'b111111111111;
		12'b001101010011: color_data = 12'b111111111111;
		12'b001101010100: color_data = 12'b000000000000;
		12'b001101010101: color_data = 12'b111111111111;
		12'b001101010110: color_data = 12'b111111111111;
		12'b001101010111: color_data = 12'b111111111111;
		12'b001101011000: color_data = 12'b111111111111;
		12'b001101011001: color_data = 12'b111111111111;
		12'b001101011010: color_data = 12'b000000000000;
		12'b001101011011: color_data = 12'b111111111111;
		12'b001101011100: color_data = 12'b111111111111;
		12'b001101011101: color_data = 12'b111111111111;
		12'b001101011110: color_data = 12'b111111111111;
		12'b001101011111: color_data = 12'b111111111111;

		12'b001101100000: color_data = 12'b111111111111;
		12'b001101100001: color_data = 12'b111111111111;
		12'b001101100010: color_data = 12'b111111111111;
		12'b001101100011: color_data = 12'b111111111111;
		12'b001101100100: color_data = 12'b111111111111;
		12'b001101100101: color_data = 12'b111111111111;
		12'b001101100110: color_data = 12'b111111111111;
		12'b001101100111: color_data = 12'b111111111111;
		12'b001101101000: color_data = 12'b111111111111;
		12'b001101101001: color_data = 12'b111111111111;
		12'b001101101010: color_data = 12'b000000000000;
		12'b001101101011: color_data = 12'b111111111111;
		12'b001101101100: color_data = 12'b111111111111;
		12'b001101101101: color_data = 12'b111111111111;
		12'b001101101110: color_data = 12'b111111111111;
		12'b001101101111: color_data = 12'b111111111111;

		12'b001101110000: color_data = 12'b111111111111;
		12'b001101110001: color_data = 12'b111111111111;
		12'b001101110010: color_data = 12'b111111111111;
		12'b001101110011: color_data = 12'b111111111111;
		12'b001101110100: color_data = 12'b111111111111;
		12'b001101110101: color_data = 12'b111111111111;
		12'b001101110110: color_data = 12'b111111111111;
		12'b001101110111: color_data = 12'b111111111111;
		12'b001101111000: color_data = 12'b111111111111;
		12'b001101111001: color_data = 12'b111111111111;
		12'b001101111010: color_data = 12'b000000000000;
		12'b001101111011: color_data = 12'b111111111111;
		12'b001101111100: color_data = 12'b111111111111;
		12'b001101111101: color_data = 12'b111111111111;
		12'b001101111110: color_data = 12'b111111111111;
		12'b001101111111: color_data = 12'b111111111111;

		12'b001110000000: color_data = 12'b111111111111;
		12'b001110000001: color_data = 12'b111111111111;
		12'b001110000010: color_data = 12'b111111111111;
		12'b001110000011: color_data = 12'b111111111111;
		12'b001110000100: color_data = 12'b111111111111;
		12'b001110000101: color_data = 12'b111111111111;
		12'b001110000110: color_data = 12'b111111111111;
		12'b001110000111: color_data = 12'b111111111111;
		12'b001110001000: color_data = 12'b111111111111;
		12'b001110001001: color_data = 12'b111111111111;
		12'b001110001010: color_data = 12'b000000000000;
		12'b001110001011: color_data = 12'b111111111111;
		12'b001110001100: color_data = 12'b111111111111;
		12'b001110001101: color_data = 12'b111111111111;
		12'b001110001110: color_data = 12'b111111111111;
		12'b001110001111: color_data = 12'b111111111111;

		12'b001110010000: color_data = 12'b111111111111;
		12'b001110010001: color_data = 12'b111111111111;
		12'b001110010010: color_data = 12'b111111111111;
		12'b001110010011: color_data = 12'b111111111111;
		12'b001110010100: color_data = 12'b000000000000;
		12'b001110010101: color_data = 12'b000000000000;
		12'b001110010110: color_data = 12'b000000000000;
		12'b001110010111: color_data = 12'b000000000000;
		12'b001110011000: color_data = 12'b000000000000;
		12'b001110011001: color_data = 12'b000000000000;
		12'b001110011010: color_data = 12'b000000000000;
		12'b001110011011: color_data = 12'b111111111111;
		12'b001110011100: color_data = 12'b111111111111;
		12'b001110011101: color_data = 12'b111111111111;
		12'b001110011110: color_data = 12'b111111111111;
		12'b001110011111: color_data = 12'b111111111111;

		12'b001110100000: color_data = 12'b111111111111;
		12'b001110100001: color_data = 12'b111111111111;
		12'b001110100010: color_data = 12'b111111111111;
		12'b001110100011: color_data = 12'b111111111111;
		12'b001110100100: color_data = 12'b111111111111;
		12'b001110100101: color_data = 12'b111111111111;
		12'b001110100110: color_data = 12'b111111111111;
		12'b001110100111: color_data = 12'b111111111111;
		12'b001110101000: color_data = 12'b111111111111;
		12'b001110101001: color_data = 12'b111111111111;
		12'b001110101010: color_data = 12'b000000000000;
		12'b001110101011: color_data = 12'b111111111111;
		12'b001110101100: color_data = 12'b111111111111;
		12'b001110101101: color_data = 12'b111111111111;
		12'b001110101110: color_data = 12'b111111111111;
		12'b001110101111: color_data = 12'b111111111111;

		12'b001110110000: color_data = 12'b111111111111;
		12'b001110110001: color_data = 12'b111111111111;
		12'b001110110010: color_data = 12'b111111111111;
		12'b001110110011: color_data = 12'b111111111111;
		12'b001110110100: color_data = 12'b111111111111;
		12'b001110110101: color_data = 12'b111111111111;
		12'b001110110110: color_data = 12'b111111111111;
		12'b001110110111: color_data = 12'b111111111111;
		12'b001110111000: color_data = 12'b111111111111;
		12'b001110111001: color_data = 12'b111111111111;
		12'b001110111010: color_data = 12'b000000000000;
		12'b001110111011: color_data = 12'b111111111111;
		12'b001110111100: color_data = 12'b111111111111;
		12'b001110111101: color_data = 12'b111111111111;
		12'b001110111110: color_data = 12'b111111111111;
		12'b001110111111: color_data = 12'b111111111111;

		12'b001111000000: color_data = 12'b111111111111;
		12'b001111000001: color_data = 12'b111111111111;
		12'b001111000010: color_data = 12'b111111111111;
		12'b001111000011: color_data = 12'b111111111111;
		12'b001111000100: color_data = 12'b111111111111;
		12'b001111000101: color_data = 12'b111111111111;
		12'b001111000110: color_data = 12'b111111111111;
		12'b001111000111: color_data = 12'b111111111111;
		12'b001111001000: color_data = 12'b111111111111;
		12'b001111001001: color_data = 12'b111111111111;
		12'b001111001010: color_data = 12'b000000000000;
		12'b001111001011: color_data = 12'b111111111111;
		12'b001111001100: color_data = 12'b111111111111;
		12'b001111001101: color_data = 12'b111111111111;
		12'b001111001110: color_data = 12'b111111111111;
		12'b001111001111: color_data = 12'b111111111111;

		12'b001111010000: color_data = 12'b111111111111;
		12'b001111010001: color_data = 12'b111111111111;
		12'b001111010010: color_data = 12'b111111111111;
		12'b001111010011: color_data = 12'b111111111111;
		12'b001111010100: color_data = 12'b000000000000;
		12'b001111010101: color_data = 12'b000000000000;
		12'b001111010110: color_data = 12'b000000000000;
		12'b001111010111: color_data = 12'b000000000000;
		12'b001111011000: color_data = 12'b000000000000;
		12'b001111011001: color_data = 12'b000000000000;
		12'b001111011010: color_data = 12'b000000000000;
		12'b001111011011: color_data = 12'b111111111111;
		12'b001111011100: color_data = 12'b111111111111;
		12'b001111011101: color_data = 12'b111111111111;
		12'b001111011110: color_data = 12'b111111111111;
		12'b001111011111: color_data = 12'b111111111111;

		12'b001111100000: color_data = 12'b111111111111;
		12'b001111100001: color_data = 12'b111111111111;
		12'b001111100010: color_data = 12'b111111111111;
		12'b001111100011: color_data = 12'b111111111111;
		12'b001111100100: color_data = 12'b111111111111;
		12'b001111100101: color_data = 12'b111111111111;
		12'b001111100110: color_data = 12'b111111111111;
		12'b001111100111: color_data = 12'b111111111111;
		12'b001111101000: color_data = 12'b111111111111;
		12'b001111101001: color_data = 12'b111111111111;
		12'b001111101010: color_data = 12'b111111111111;
		12'b001111101011: color_data = 12'b111111111111;
		12'b001111101100: color_data = 12'b111111111111;
		12'b001111101101: color_data = 12'b111111111111;
		12'b001111101110: color_data = 12'b111111111111;
		12'b001111101111: color_data = 12'b111111111111;

		12'b001111110000: color_data = 12'b111111111111;
		12'b001111110001: color_data = 12'b111111111111;
		12'b001111110010: color_data = 12'b111111111111;
		12'b001111110011: color_data = 12'b111111111111;
		12'b001111110100: color_data = 12'b111111111111;
		12'b001111110101: color_data = 12'b111111111111;
		12'b001111110110: color_data = 12'b111111111111;
		12'b001111110111: color_data = 12'b111111111111;
		12'b001111111000: color_data = 12'b111111111111;
		12'b001111111001: color_data = 12'b111111111111;
		12'b001111111010: color_data = 12'b111111111111;
		12'b001111111011: color_data = 12'b111111111111;
		12'b001111111100: color_data = 12'b111111111111;
		12'b001111111101: color_data = 12'b111111111111;
		12'b001111111110: color_data = 12'b111111111111;
		12'b001111111111: color_data = 12'b111111111111;

		12'b010000000000: color_data = 12'b111111111111;
		12'b010000000001: color_data = 12'b111111111111;
		12'b010000000010: color_data = 12'b111111111111;
		12'b010000000011: color_data = 12'b111111111111;
		12'b010000000100: color_data = 12'b111111111111;
		12'b010000000101: color_data = 12'b111111111111;
		12'b010000000110: color_data = 12'b111111111111;
		12'b010000000111: color_data = 12'b111111111111;
		12'b010000001000: color_data = 12'b111111111111;
		12'b010000001001: color_data = 12'b111111111111;
		12'b010000001010: color_data = 12'b111111111111;
		12'b010000001011: color_data = 12'b111111111111;
		12'b010000001100: color_data = 12'b111111111111;
		12'b010000001101: color_data = 12'b111111111111;
		12'b010000001110: color_data = 12'b111111111111;
		12'b010000001111: color_data = 12'b111111111111;

		12'b010000010000: color_data = 12'b111111111111;
		12'b010000010001: color_data = 12'b111111111111;
		12'b010000010010: color_data = 12'b111111111111;
		12'b010000010011: color_data = 12'b111111111111;
		12'b010000010100: color_data = 12'b000000000000;
		12'b010000010101: color_data = 12'b111111111111;
		12'b010000010110: color_data = 12'b111111111111;
		12'b010000010111: color_data = 12'b111111111111;
		12'b010000011000: color_data = 12'b111111111111;
		12'b010000011001: color_data = 12'b111111111111;
		12'b010000011010: color_data = 12'b000000000000;
		12'b010000011011: color_data = 12'b111111111111;
		12'b010000011100: color_data = 12'b111111111111;
		12'b010000011101: color_data = 12'b111111111111;
		12'b010000011110: color_data = 12'b111111111111;
		12'b010000011111: color_data = 12'b111111111111;

		12'b010000100000: color_data = 12'b111111111111;
		12'b010000100001: color_data = 12'b111111111111;
		12'b010000100010: color_data = 12'b111111111111;
		12'b010000100011: color_data = 12'b111111111111;
		12'b010000100100: color_data = 12'b000000000000;
		12'b010000100101: color_data = 12'b111111111111;
		12'b010000100110: color_data = 12'b111111111111;
		12'b010000100111: color_data = 12'b111111111111;
		12'b010000101000: color_data = 12'b111111111111;
		12'b010000101001: color_data = 12'b111111111111;
		12'b010000101010: color_data = 12'b000000000000;
		12'b010000101011: color_data = 12'b111111111111;
		12'b010000101100: color_data = 12'b111111111111;
		12'b010000101101: color_data = 12'b111111111111;
		12'b010000101110: color_data = 12'b111111111111;
		12'b010000101111: color_data = 12'b111111111111;

		12'b010000110000: color_data = 12'b111111111111;
		12'b010000110001: color_data = 12'b111111111111;
		12'b010000110010: color_data = 12'b111111111111;
		12'b010000110011: color_data = 12'b111111111111;
		12'b010000110100: color_data = 12'b000000000000;
		12'b010000110101: color_data = 12'b111111111111;
		12'b010000110110: color_data = 12'b111111111111;
		12'b010000110111: color_data = 12'b111111111111;
		12'b010000111000: color_data = 12'b111111111111;
		12'b010000111001: color_data = 12'b111111111111;
		12'b010000111010: color_data = 12'b000000000000;
		12'b010000111011: color_data = 12'b111111111111;
		12'b010000111100: color_data = 12'b111111111111;
		12'b010000111101: color_data = 12'b111111111111;
		12'b010000111110: color_data = 12'b111111111111;
		12'b010000111111: color_data = 12'b111111111111;

		12'b010001000000: color_data = 12'b111111111111;
		12'b010001000001: color_data = 12'b111111111111;
		12'b010001000010: color_data = 12'b111111111111;
		12'b010001000011: color_data = 12'b111111111111;
		12'b010001000100: color_data = 12'b000000000000;
		12'b010001000101: color_data = 12'b111111111111;
		12'b010001000110: color_data = 12'b111111111111;
		12'b010001000111: color_data = 12'b111111111111;
		12'b010001001000: color_data = 12'b111111111111;
		12'b010001001001: color_data = 12'b111111111111;
		12'b010001001010: color_data = 12'b000000000000;
		12'b010001001011: color_data = 12'b111111111111;
		12'b010001001100: color_data = 12'b111111111111;
		12'b010001001101: color_data = 12'b111111111111;
		12'b010001001110: color_data = 12'b111111111111;
		12'b010001001111: color_data = 12'b111111111111;

		12'b010001010000: color_data = 12'b111111111111;
		12'b010001010001: color_data = 12'b111111111111;
		12'b010001010010: color_data = 12'b111111111111;
		12'b010001010011: color_data = 12'b111111111111;
		12'b010001010100: color_data = 12'b000000000000;
		12'b010001010101: color_data = 12'b111111111111;
		12'b010001010110: color_data = 12'b111111111111;
		12'b010001010111: color_data = 12'b111111111111;
		12'b010001011000: color_data = 12'b111111111111;
		12'b010001011001: color_data = 12'b111111111111;
		12'b010001011010: color_data = 12'b000000000000;
		12'b010001011011: color_data = 12'b111111111111;
		12'b010001011100: color_data = 12'b111111111111;
		12'b010001011101: color_data = 12'b111111111111;
		12'b010001011110: color_data = 12'b111111111111;
		12'b010001011111: color_data = 12'b111111111111;

		12'b010001100000: color_data = 12'b111111111111;
		12'b010001100001: color_data = 12'b111111111111;
		12'b010001100010: color_data = 12'b111111111111;
		12'b010001100011: color_data = 12'b111111111111;
		12'b010001100100: color_data = 12'b000000000000;
		12'b010001100101: color_data = 12'b111111111111;
		12'b010001100110: color_data = 12'b111111111111;
		12'b010001100111: color_data = 12'b111111111111;
		12'b010001101000: color_data = 12'b111111111111;
		12'b010001101001: color_data = 12'b111111111111;
		12'b010001101010: color_data = 12'b000000000000;
		12'b010001101011: color_data = 12'b111111111111;
		12'b010001101100: color_data = 12'b111111111111;
		12'b010001101101: color_data = 12'b111111111111;
		12'b010001101110: color_data = 12'b111111111111;
		12'b010001101111: color_data = 12'b111111111111;

		12'b010001110000: color_data = 12'b111111111111;
		12'b010001110001: color_data = 12'b111111111111;
		12'b010001110010: color_data = 12'b111111111111;
		12'b010001110011: color_data = 12'b111111111111;
		12'b010001110100: color_data = 12'b000000000000;
		12'b010001110101: color_data = 12'b000000000000;
		12'b010001110110: color_data = 12'b000000000000;
		12'b010001110111: color_data = 12'b000000000000;
		12'b010001111000: color_data = 12'b000000000000;
		12'b010001111001: color_data = 12'b000000000000;
		12'b010001111010: color_data = 12'b000000000000;
		12'b010001111011: color_data = 12'b111111111111;
		12'b010001111100: color_data = 12'b111111111111;
		12'b010001111101: color_data = 12'b111111111111;
		12'b010001111110: color_data = 12'b111111111111;
		12'b010001111111: color_data = 12'b111111111111;

		12'b010010000000: color_data = 12'b111111111111;
		12'b010010000001: color_data = 12'b111111111111;
		12'b010010000010: color_data = 12'b111111111111;
		12'b010010000011: color_data = 12'b111111111111;
		12'b010010000100: color_data = 12'b111111111111;
		12'b010010000101: color_data = 12'b111111111111;
		12'b010010000110: color_data = 12'b111111111111;
		12'b010010000111: color_data = 12'b111111111111;
		12'b010010001000: color_data = 12'b111111111111;
		12'b010010001001: color_data = 12'b111111111111;
		12'b010010001010: color_data = 12'b000000000000;
		12'b010010001011: color_data = 12'b111111111111;
		12'b010010001100: color_data = 12'b111111111111;
		12'b010010001101: color_data = 12'b111111111111;
		12'b010010001110: color_data = 12'b111111111111;
		12'b010010001111: color_data = 12'b111111111111;

		12'b010010010000: color_data = 12'b111111111111;
		12'b010010010001: color_data = 12'b111111111111;
		12'b010010010010: color_data = 12'b111111111111;
		12'b010010010011: color_data = 12'b111111111111;
		12'b010010010100: color_data = 12'b111111111111;
		12'b010010010101: color_data = 12'b111111111111;
		12'b010010010110: color_data = 12'b111111111111;
		12'b010010010111: color_data = 12'b111111111111;
		12'b010010011000: color_data = 12'b111111111111;
		12'b010010011001: color_data = 12'b111111111111;
		12'b010010011010: color_data = 12'b000000000000;
		12'b010010011011: color_data = 12'b111111111111;
		12'b010010011100: color_data = 12'b111111111111;
		12'b010010011101: color_data = 12'b111111111111;
		12'b010010011110: color_data = 12'b111111111111;
		12'b010010011111: color_data = 12'b111111111111;

		12'b010010100000: color_data = 12'b111111111111;
		12'b010010100001: color_data = 12'b111111111111;
		12'b010010100010: color_data = 12'b111111111111;
		12'b010010100011: color_data = 12'b111111111111;
		12'b010010100100: color_data = 12'b111111111111;
		12'b010010100101: color_data = 12'b111111111111;
		12'b010010100110: color_data = 12'b111111111111;
		12'b010010100111: color_data = 12'b111111111111;
		12'b010010101000: color_data = 12'b111111111111;
		12'b010010101001: color_data = 12'b111111111111;
		12'b010010101010: color_data = 12'b000000000000;
		12'b010010101011: color_data = 12'b111111111111;
		12'b010010101100: color_data = 12'b111111111111;
		12'b010010101101: color_data = 12'b111111111111;
		12'b010010101110: color_data = 12'b111111111111;
		12'b010010101111: color_data = 12'b111111111111;

		12'b010010110000: color_data = 12'b111111111111;
		12'b010010110001: color_data = 12'b111111111111;
		12'b010010110010: color_data = 12'b111111111111;
		12'b010010110011: color_data = 12'b111111111111;
		12'b010010110100: color_data = 12'b111111111111;
		12'b010010110101: color_data = 12'b111111111111;
		12'b010010110110: color_data = 12'b111111111111;
		12'b010010110111: color_data = 12'b111111111111;
		12'b010010111000: color_data = 12'b111111111111;
		12'b010010111001: color_data = 12'b111111111111;
		12'b010010111010: color_data = 12'b000000000000;
		12'b010010111011: color_data = 12'b111111111111;
		12'b010010111100: color_data = 12'b111111111111;
		12'b010010111101: color_data = 12'b111111111111;
		12'b010010111110: color_data = 12'b111111111111;
		12'b010010111111: color_data = 12'b111111111111;

		12'b010011000000: color_data = 12'b111111111111;
		12'b010011000001: color_data = 12'b111111111111;
		12'b010011000010: color_data = 12'b111111111111;
		12'b010011000011: color_data = 12'b111111111111;
		12'b010011000100: color_data = 12'b111111111111;
		12'b010011000101: color_data = 12'b111111111111;
		12'b010011000110: color_data = 12'b111111111111;
		12'b010011000111: color_data = 12'b111111111111;
		12'b010011001000: color_data = 12'b111111111111;
		12'b010011001001: color_data = 12'b111111111111;
		12'b010011001010: color_data = 12'b000000000000;
		12'b010011001011: color_data = 12'b111111111111;
		12'b010011001100: color_data = 12'b111111111111;
		12'b010011001101: color_data = 12'b111111111111;
		12'b010011001110: color_data = 12'b111111111111;
		12'b010011001111: color_data = 12'b111111111111;

		12'b010011010000: color_data = 12'b111111111111;
		12'b010011010001: color_data = 12'b111111111111;
		12'b010011010010: color_data = 12'b111111111111;
		12'b010011010011: color_data = 12'b111111111111;
		12'b010011010100: color_data = 12'b111111111111;
		12'b010011010101: color_data = 12'b111111111111;
		12'b010011010110: color_data = 12'b111111111111;
		12'b010011010111: color_data = 12'b111111111111;
		12'b010011011000: color_data = 12'b111111111111;
		12'b010011011001: color_data = 12'b111111111111;
		12'b010011011010: color_data = 12'b000000000000;
		12'b010011011011: color_data = 12'b111111111111;
		12'b010011011100: color_data = 12'b111111111111;
		12'b010011011101: color_data = 12'b111111111111;
		12'b010011011110: color_data = 12'b111111111111;
		12'b010011011111: color_data = 12'b111111111111;

		12'b010011100000: color_data = 12'b111111111111;
		12'b010011100001: color_data = 12'b111111111111;
		12'b010011100010: color_data = 12'b111111111111;
		12'b010011100011: color_data = 12'b111111111111;
		12'b010011100100: color_data = 12'b111111111111;
		12'b010011100101: color_data = 12'b111111111111;
		12'b010011100110: color_data = 12'b111111111111;
		12'b010011100111: color_data = 12'b111111111111;
		12'b010011101000: color_data = 12'b111111111111;
		12'b010011101001: color_data = 12'b111111111111;
		12'b010011101010: color_data = 12'b111111111111;
		12'b010011101011: color_data = 12'b111111111111;
		12'b010011101100: color_data = 12'b111111111111;
		12'b010011101101: color_data = 12'b111111111111;
		12'b010011101110: color_data = 12'b111111111111;
		12'b010011101111: color_data = 12'b111111111111;

		12'b010011110000: color_data = 12'b111111111111;
		12'b010011110001: color_data = 12'b111111111111;
		12'b010011110010: color_data = 12'b111111111111;
		12'b010011110011: color_data = 12'b111111111111;
		12'b010011110100: color_data = 12'b111111111111;
		12'b010011110101: color_data = 12'b111111111111;
		12'b010011110110: color_data = 12'b111111111111;
		12'b010011110111: color_data = 12'b111111111111;
		12'b010011111000: color_data = 12'b111111111111;
		12'b010011111001: color_data = 12'b111111111111;
		12'b010011111010: color_data = 12'b111111111111;
		12'b010011111011: color_data = 12'b111111111111;
		12'b010011111100: color_data = 12'b111111111111;
		12'b010011111101: color_data = 12'b111111111111;
		12'b010011111110: color_data = 12'b111111111111;
		12'b010011111111: color_data = 12'b111111111111;

		12'b010100000000: color_data = 12'b111111111111;
		12'b010100000001: color_data = 12'b111111111111;
		12'b010100000010: color_data = 12'b111111111111;
		12'b010100000011: color_data = 12'b111111111111;
		12'b010100000100: color_data = 12'b111111111111;
		12'b010100000101: color_data = 12'b111111111111;
		12'b010100000110: color_data = 12'b111111111111;
		12'b010100000111: color_data = 12'b111111111111;
		12'b010100001000: color_data = 12'b111111111111;
		12'b010100001001: color_data = 12'b111111111111;
		12'b010100001010: color_data = 12'b111111111111;
		12'b010100001011: color_data = 12'b111111111111;
		12'b010100001100: color_data = 12'b111111111111;
		12'b010100001101: color_data = 12'b111111111111;
		12'b010100001110: color_data = 12'b111111111111;
		12'b010100001111: color_data = 12'b111111111111;

		12'b010100010000: color_data = 12'b111111111111;
		12'b010100010001: color_data = 12'b111111111111;
		12'b010100010010: color_data = 12'b111111111111;
		12'b010100010011: color_data = 12'b111111111111;
		12'b010100010100: color_data = 12'b000000000000;
		12'b010100010101: color_data = 12'b000000000000;
		12'b010100010110: color_data = 12'b000000000000;
		12'b010100010111: color_data = 12'b000000000000;
		12'b010100011000: color_data = 12'b000000000000;
		12'b010100011001: color_data = 12'b000000000000;
		12'b010100011010: color_data = 12'b000000000000;
		12'b010100011011: color_data = 12'b111111111111;
		12'b010100011100: color_data = 12'b111111111111;
		12'b010100011101: color_data = 12'b111111111111;
		12'b010100011110: color_data = 12'b111111111111;
		12'b010100011111: color_data = 12'b111111111111;

		12'b010100100000: color_data = 12'b111111111111;
		12'b010100100001: color_data = 12'b111111111111;
		12'b010100100010: color_data = 12'b111111111111;
		12'b010100100011: color_data = 12'b111111111111;
		12'b010100100100: color_data = 12'b000000000000;
		12'b010100100101: color_data = 12'b111111111111;
		12'b010100100110: color_data = 12'b111111111111;
		12'b010100100111: color_data = 12'b111111111111;
		12'b010100101000: color_data = 12'b111111111111;
		12'b010100101001: color_data = 12'b111111111111;
		12'b010100101010: color_data = 12'b111111111111;
		12'b010100101011: color_data = 12'b111111111111;
		12'b010100101100: color_data = 12'b111111111111;
		12'b010100101101: color_data = 12'b111111111111;
		12'b010100101110: color_data = 12'b111111111111;
		12'b010100101111: color_data = 12'b111111111111;

		12'b010100110000: color_data = 12'b111111111111;
		12'b010100110001: color_data = 12'b111111111111;
		12'b010100110010: color_data = 12'b111111111111;
		12'b010100110011: color_data = 12'b111111111111;
		12'b010100110100: color_data = 12'b000000000000;
		12'b010100110101: color_data = 12'b111111111111;
		12'b010100110110: color_data = 12'b111111111111;
		12'b010100110111: color_data = 12'b111111111111;
		12'b010100111000: color_data = 12'b111111111111;
		12'b010100111001: color_data = 12'b111111111111;
		12'b010100111010: color_data = 12'b111111111111;
		12'b010100111011: color_data = 12'b111111111111;
		12'b010100111100: color_data = 12'b111111111111;
		12'b010100111101: color_data = 12'b111111111111;
		12'b010100111110: color_data = 12'b111111111111;
		12'b010100111111: color_data = 12'b111111111111;

		12'b010101000000: color_data = 12'b111111111111;
		12'b010101000001: color_data = 12'b111111111111;
		12'b010101000010: color_data = 12'b111111111111;
		12'b010101000011: color_data = 12'b111111111111;
		12'b010101000100: color_data = 12'b000000000000;
		12'b010101000101: color_data = 12'b111111111111;
		12'b010101000110: color_data = 12'b111111111111;
		12'b010101000111: color_data = 12'b111111111111;
		12'b010101001000: color_data = 12'b111111111111;
		12'b010101001001: color_data = 12'b111111111111;
		12'b010101001010: color_data = 12'b111111111111;
		12'b010101001011: color_data = 12'b111111111111;
		12'b010101001100: color_data = 12'b111111111111;
		12'b010101001101: color_data = 12'b111111111111;
		12'b010101001110: color_data = 12'b111111111111;
		12'b010101001111: color_data = 12'b111111111111;

		12'b010101010000: color_data = 12'b111111111111;
		12'b010101010001: color_data = 12'b111111111111;
		12'b010101010010: color_data = 12'b111111111111;
		12'b010101010011: color_data = 12'b111111111111;
		12'b010101010100: color_data = 12'b000000000000;
		12'b010101010101: color_data = 12'b111111111111;
		12'b010101010110: color_data = 12'b111111111111;
		12'b010101010111: color_data = 12'b111111111111;
		12'b010101011000: color_data = 12'b111111111111;
		12'b010101011001: color_data = 12'b111111111111;
		12'b010101011010: color_data = 12'b111111111111;
		12'b010101011011: color_data = 12'b111111111111;
		12'b010101011100: color_data = 12'b111111111111;
		12'b010101011101: color_data = 12'b111111111111;
		12'b010101011110: color_data = 12'b111111111111;
		12'b010101011111: color_data = 12'b111111111111;

		12'b010101100000: color_data = 12'b111111111111;
		12'b010101100001: color_data = 12'b111111111111;
		12'b010101100010: color_data = 12'b111111111111;
		12'b010101100011: color_data = 12'b111111111111;
		12'b010101100100: color_data = 12'b000000000000;
		12'b010101100101: color_data = 12'b111111111111;
		12'b010101100110: color_data = 12'b111111111111;
		12'b010101100111: color_data = 12'b111111111111;
		12'b010101101000: color_data = 12'b111111111111;
		12'b010101101001: color_data = 12'b111111111111;
		12'b010101101010: color_data = 12'b111111111111;
		12'b010101101011: color_data = 12'b111111111111;
		12'b010101101100: color_data = 12'b111111111111;
		12'b010101101101: color_data = 12'b111111111111;
		12'b010101101110: color_data = 12'b111111111111;
		12'b010101101111: color_data = 12'b111111111111;

		12'b010101110000: color_data = 12'b111111111111;
		12'b010101110001: color_data = 12'b111111111111;
		12'b010101110010: color_data = 12'b111111111111;
		12'b010101110011: color_data = 12'b111111111111;
		12'b010101110100: color_data = 12'b000000000000;
		12'b010101110101: color_data = 12'b111111111111;
		12'b010101110110: color_data = 12'b111111111111;
		12'b010101110111: color_data = 12'b111111111111;
		12'b010101111000: color_data = 12'b111111111111;
		12'b010101111001: color_data = 12'b111111111111;
		12'b010101111010: color_data = 12'b111111111111;
		12'b010101111011: color_data = 12'b111111111111;
		12'b010101111100: color_data = 12'b111111111111;
		12'b010101111101: color_data = 12'b111111111111;
		12'b010101111110: color_data = 12'b111111111111;
		12'b010101111111: color_data = 12'b111111111111;

		12'b010110000000: color_data = 12'b111111111111;
		12'b010110000001: color_data = 12'b111111111111;
		12'b010110000010: color_data = 12'b111111111111;
		12'b010110000011: color_data = 12'b111111111111;
		12'b010110000100: color_data = 12'b000000000000;
		12'b010110000101: color_data = 12'b000000000000;
		12'b010110000110: color_data = 12'b000000000000;
		12'b010110000111: color_data = 12'b000000000000;
		12'b010110001000: color_data = 12'b000000000000;
		12'b010110001001: color_data = 12'b000000000000;
		12'b010110001010: color_data = 12'b000000000000;
		12'b010110001011: color_data = 12'b111111111111;
		12'b010110001100: color_data = 12'b111111111111;
		12'b010110001101: color_data = 12'b111111111111;
		12'b010110001110: color_data = 12'b111111111111;
		12'b010110001111: color_data = 12'b111111111111;

		12'b010110010000: color_data = 12'b111111111111;
		12'b010110010001: color_data = 12'b111111111111;
		12'b010110010010: color_data = 12'b111111111111;
		12'b010110010011: color_data = 12'b111111111111;
		12'b010110010100: color_data = 12'b111111111111;
		12'b010110010101: color_data = 12'b111111111111;
		12'b010110010110: color_data = 12'b111111111111;
		12'b010110010111: color_data = 12'b111111111111;
		12'b010110011000: color_data = 12'b111111111111;
		12'b010110011001: color_data = 12'b111111111111;
		12'b010110011010: color_data = 12'b000000000000;
		12'b010110011011: color_data = 12'b111111111111;
		12'b010110011100: color_data = 12'b111111111111;
		12'b010110011101: color_data = 12'b111111111111;
		12'b010110011110: color_data = 12'b111111111111;
		12'b010110011111: color_data = 12'b111111111111;

		12'b010110100000: color_data = 12'b111111111111;
		12'b010110100001: color_data = 12'b111111111111;
		12'b010110100010: color_data = 12'b111111111111;
		12'b010110100011: color_data = 12'b111111111111;
		12'b010110100100: color_data = 12'b111111111111;
		12'b010110100101: color_data = 12'b111111111111;
		12'b010110100110: color_data = 12'b111111111111;
		12'b010110100111: color_data = 12'b111111111111;
		12'b010110101000: color_data = 12'b111111111111;
		12'b010110101001: color_data = 12'b111111111111;
		12'b010110101010: color_data = 12'b000000000000;
		12'b010110101011: color_data = 12'b111111111111;
		12'b010110101100: color_data = 12'b111111111111;
		12'b010110101101: color_data = 12'b111111111111;
		12'b010110101110: color_data = 12'b111111111111;
		12'b010110101111: color_data = 12'b111111111111;

		12'b010110110000: color_data = 12'b111111111111;
		12'b010110110001: color_data = 12'b111111111111;
		12'b010110110010: color_data = 12'b111111111111;
		12'b010110110011: color_data = 12'b111111111111;
		12'b010110110100: color_data = 12'b111111111111;
		12'b010110110101: color_data = 12'b111111111111;
		12'b010110110110: color_data = 12'b111111111111;
		12'b010110110111: color_data = 12'b111111111111;
		12'b010110111000: color_data = 12'b111111111111;
		12'b010110111001: color_data = 12'b111111111111;
		12'b010110111010: color_data = 12'b000000000000;
		12'b010110111011: color_data = 12'b111111111111;
		12'b010110111100: color_data = 12'b111111111111;
		12'b010110111101: color_data = 12'b111111111111;
		12'b010110111110: color_data = 12'b111111111111;
		12'b010110111111: color_data = 12'b111111111111;

		12'b010111000000: color_data = 12'b111111111111;
		12'b010111000001: color_data = 12'b111111111111;
		12'b010111000010: color_data = 12'b111111111111;
		12'b010111000011: color_data = 12'b111111111111;
		12'b010111000100: color_data = 12'b111111111111;
		12'b010111000101: color_data = 12'b111111111111;
		12'b010111000110: color_data = 12'b111111111111;
		12'b010111000111: color_data = 12'b111111111111;
		12'b010111001000: color_data = 12'b111111111111;
		12'b010111001001: color_data = 12'b111111111111;
		12'b010111001010: color_data = 12'b000000000000;
		12'b010111001011: color_data = 12'b111111111111;
		12'b010111001100: color_data = 12'b111111111111;
		12'b010111001101: color_data = 12'b111111111111;
		12'b010111001110: color_data = 12'b111111111111;
		12'b010111001111: color_data = 12'b111111111111;

		12'b010111010000: color_data = 12'b111111111111;
		12'b010111010001: color_data = 12'b111111111111;
		12'b010111010010: color_data = 12'b111111111111;
		12'b010111010011: color_data = 12'b111111111111;
		12'b010111010100: color_data = 12'b000000000000;
		12'b010111010101: color_data = 12'b000000000000;
		12'b010111010110: color_data = 12'b000000000000;
		12'b010111010111: color_data = 12'b000000000000;
		12'b010111011000: color_data = 12'b000000000000;
		12'b010111011001: color_data = 12'b000000000000;
		12'b010111011010: color_data = 12'b000000000000;
		12'b010111011011: color_data = 12'b111111111111;
		12'b010111011100: color_data = 12'b111111111111;
		12'b010111011101: color_data = 12'b111111111111;
		12'b010111011110: color_data = 12'b111111111111;
		12'b010111011111: color_data = 12'b111111111111;

		12'b010111100000: color_data = 12'b111111111111;
		12'b010111100001: color_data = 12'b111111111111;
		12'b010111100010: color_data = 12'b111111111111;
		12'b010111100011: color_data = 12'b111111111111;
		12'b010111100100: color_data = 12'b111111111111;
		12'b010111100101: color_data = 12'b111111111111;
		12'b010111100110: color_data = 12'b111111111111;
		12'b010111100111: color_data = 12'b111111111111;
		12'b010111101000: color_data = 12'b111111111111;
		12'b010111101001: color_data = 12'b111111111111;
		12'b010111101010: color_data = 12'b111111111111;
		12'b010111101011: color_data = 12'b111111111111;
		12'b010111101100: color_data = 12'b111111111111;
		12'b010111101101: color_data = 12'b111111111111;
		12'b010111101110: color_data = 12'b111111111111;
		12'b010111101111: color_data = 12'b111111111111;

		12'b010111110000: color_data = 12'b111111111111;
		12'b010111110001: color_data = 12'b111111111111;
		12'b010111110010: color_data = 12'b111111111111;
		12'b010111110011: color_data = 12'b111111111111;
		12'b010111110100: color_data = 12'b111111111111;
		12'b010111110101: color_data = 12'b111111111111;
		12'b010111110110: color_data = 12'b111111111111;
		12'b010111110111: color_data = 12'b111111111111;
		12'b010111111000: color_data = 12'b111111111111;
		12'b010111111001: color_data = 12'b111111111111;
		12'b010111111010: color_data = 12'b111111111111;
		12'b010111111011: color_data = 12'b111111111111;
		12'b010111111100: color_data = 12'b111111111111;
		12'b010111111101: color_data = 12'b111111111111;
		12'b010111111110: color_data = 12'b111111111111;
		12'b010111111111: color_data = 12'b111111111111;

		12'b011000000000: color_data = 12'b111111111111;
		12'b011000000001: color_data = 12'b111111111111;
		12'b011000000010: color_data = 12'b111111111111;
		12'b011000000011: color_data = 12'b111111111111;
		12'b011000000100: color_data = 12'b111111111111;
		12'b011000000101: color_data = 12'b111111111111;
		12'b011000000110: color_data = 12'b111111111111;
		12'b011000000111: color_data = 12'b111111111111;
		12'b011000001000: color_data = 12'b111111111111;
		12'b011000001001: color_data = 12'b111111111111;
		12'b011000001010: color_data = 12'b111111111111;
		12'b011000001011: color_data = 12'b111111111111;
		12'b011000001100: color_data = 12'b111111111111;
		12'b011000001101: color_data = 12'b111111111111;
		12'b011000001110: color_data = 12'b111111111111;
		12'b011000001111: color_data = 12'b111111111111;

		12'b011000010000: color_data = 12'b111111111111;
		12'b011000010001: color_data = 12'b111111111111;
		12'b011000010010: color_data = 12'b111111111111;
		12'b011000010011: color_data = 12'b111111111111;
		12'b011000010100: color_data = 12'b000000000000;
		12'b011000010101: color_data = 12'b000000000000;
		12'b011000010110: color_data = 12'b000000000000;
		12'b011000010111: color_data = 12'b000000000000;
		12'b011000011000: color_data = 12'b000000000000;
		12'b011000011001: color_data = 12'b000000000000;
		12'b011000011010: color_data = 12'b000000000000;
		12'b011000011011: color_data = 12'b111111111111;
		12'b011000011100: color_data = 12'b111111111111;
		12'b011000011101: color_data = 12'b111111111111;
		12'b011000011110: color_data = 12'b111111111111;
		12'b011000011111: color_data = 12'b111111111111;

		12'b011000100000: color_data = 12'b111111111111;
		12'b011000100001: color_data = 12'b111111111111;
		12'b011000100010: color_data = 12'b111111111111;
		12'b011000100011: color_data = 12'b111111111111;
		12'b011000100100: color_data = 12'b000000000000;
		12'b011000100101: color_data = 12'b111111111111;
		12'b011000100110: color_data = 12'b111111111111;
		12'b011000100111: color_data = 12'b111111111111;
		12'b011000101000: color_data = 12'b111111111111;
		12'b011000101001: color_data = 12'b111111111111;
		12'b011000101010: color_data = 12'b000000000000;
		12'b011000101011: color_data = 12'b111111111111;
		12'b011000101100: color_data = 12'b111111111111;
		12'b011000101101: color_data = 12'b111111111111;
		12'b011000101110: color_data = 12'b111111111111;
		12'b011000101111: color_data = 12'b111111111111;

		12'b011000110000: color_data = 12'b111111111111;
		12'b011000110001: color_data = 12'b111111111111;
		12'b011000110010: color_data = 12'b111111111111;
		12'b011000110011: color_data = 12'b111111111111;
		12'b011000110100: color_data = 12'b000000000000;
		12'b011000110101: color_data = 12'b111111111111;
		12'b011000110110: color_data = 12'b111111111111;
		12'b011000110111: color_data = 12'b111111111111;
		12'b011000111000: color_data = 12'b111111111111;
		12'b011000111001: color_data = 12'b111111111111;
		12'b011000111010: color_data = 12'b000000000000;
		12'b011000111011: color_data = 12'b111111111111;
		12'b011000111100: color_data = 12'b111111111111;
		12'b011000111101: color_data = 12'b111111111111;
		12'b011000111110: color_data = 12'b111111111111;
		12'b011000111111: color_data = 12'b111111111111;

		12'b011001000000: color_data = 12'b111111111111;
		12'b011001000001: color_data = 12'b111111111111;
		12'b011001000010: color_data = 12'b111111111111;
		12'b011001000011: color_data = 12'b111111111111;
		12'b011001000100: color_data = 12'b000000000000;
		12'b011001000101: color_data = 12'b111111111111;
		12'b011001000110: color_data = 12'b111111111111;
		12'b011001000111: color_data = 12'b111111111111;
		12'b011001001000: color_data = 12'b111111111111;
		12'b011001001001: color_data = 12'b111111111111;
		12'b011001001010: color_data = 12'b111111111111;
		12'b011001001011: color_data = 12'b111111111111;
		12'b011001001100: color_data = 12'b111111111111;
		12'b011001001101: color_data = 12'b111111111111;
		12'b011001001110: color_data = 12'b111111111111;
		12'b011001001111: color_data = 12'b111111111111;

		12'b011001010000: color_data = 12'b111111111111;
		12'b011001010001: color_data = 12'b111111111111;
		12'b011001010010: color_data = 12'b111111111111;
		12'b011001010011: color_data = 12'b111111111111;
		12'b011001010100: color_data = 12'b000000000000;
		12'b011001010101: color_data = 12'b111111111111;
		12'b011001010110: color_data = 12'b111111111111;
		12'b011001010111: color_data = 12'b111111111111;
		12'b011001011000: color_data = 12'b111111111111;
		12'b011001011001: color_data = 12'b111111111111;
		12'b011001011010: color_data = 12'b111111111111;
		12'b011001011011: color_data = 12'b111111111111;
		12'b011001011100: color_data = 12'b111111111111;
		12'b011001011101: color_data = 12'b111111111111;
		12'b011001011110: color_data = 12'b111111111111;
		12'b011001011111: color_data = 12'b111111111111;

		12'b011001100000: color_data = 12'b111111111111;
		12'b011001100001: color_data = 12'b111111111111;
		12'b011001100010: color_data = 12'b111111111111;
		12'b011001100011: color_data = 12'b111111111111;
		12'b011001100100: color_data = 12'b000000000000;
		12'b011001100101: color_data = 12'b111111111111;
		12'b011001100110: color_data = 12'b111111111111;
		12'b011001100111: color_data = 12'b111111111111;
		12'b011001101000: color_data = 12'b111111111111;
		12'b011001101001: color_data = 12'b111111111111;
		12'b011001101010: color_data = 12'b111111111111;
		12'b011001101011: color_data = 12'b111111111111;
		12'b011001101100: color_data = 12'b111111111111;
		12'b011001101101: color_data = 12'b111111111111;
		12'b011001101110: color_data = 12'b111111111111;
		12'b011001101111: color_data = 12'b111111111111;

		12'b011001110000: color_data = 12'b111111111111;
		12'b011001110001: color_data = 12'b111111111111;
		12'b011001110010: color_data = 12'b111111111111;
		12'b011001110011: color_data = 12'b111111111111;
		12'b011001110100: color_data = 12'b000000000000;
		12'b011001110101: color_data = 12'b111111111111;
		12'b011001110110: color_data = 12'b111111111111;
		12'b011001110111: color_data = 12'b111111111111;
		12'b011001111000: color_data = 12'b111111111111;
		12'b011001111001: color_data = 12'b111111111111;
		12'b011001111010: color_data = 12'b111111111111;
		12'b011001111011: color_data = 12'b111111111111;
		12'b011001111100: color_data = 12'b111111111111;
		12'b011001111101: color_data = 12'b111111111111;
		12'b011001111110: color_data = 12'b111111111111;
		12'b011001111111: color_data = 12'b111111111111;

		12'b011010000000: color_data = 12'b111111111111;
		12'b011010000001: color_data = 12'b111111111111;
		12'b011010000010: color_data = 12'b111111111111;
		12'b011010000011: color_data = 12'b111111111111;
		12'b011010000100: color_data = 12'b000000000000;
		12'b011010000101: color_data = 12'b000000000000;
		12'b011010000110: color_data = 12'b000000000000;
		12'b011010000111: color_data = 12'b000000000000;
		12'b011010001000: color_data = 12'b000000000000;
		12'b011010001001: color_data = 12'b000000000000;
		12'b011010001010: color_data = 12'b000000000000;
		12'b011010001011: color_data = 12'b111111111111;
		12'b011010001100: color_data = 12'b111111111111;
		12'b011010001101: color_data = 12'b111111111111;
		12'b011010001110: color_data = 12'b111111111111;
		12'b011010001111: color_data = 12'b111111111111;

		12'b011010010000: color_data = 12'b111111111111;
		12'b011010010001: color_data = 12'b111111111111;
		12'b011010010010: color_data = 12'b111111111111;
		12'b011010010011: color_data = 12'b111111111111;
		12'b011010010100: color_data = 12'b000000000000;
		12'b011010010101: color_data = 12'b111111111111;
		12'b011010010110: color_data = 12'b111111111111;
		12'b011010010111: color_data = 12'b111111111111;
		12'b011010011000: color_data = 12'b111111111111;
		12'b011010011001: color_data = 12'b111111111111;
		12'b011010011010: color_data = 12'b000000000000;
		12'b011010011011: color_data = 12'b111111111111;
		12'b011010011100: color_data = 12'b111111111111;
		12'b011010011101: color_data = 12'b111111111111;
		12'b011010011110: color_data = 12'b111111111111;
		12'b011010011111: color_data = 12'b111111111111;

		12'b011010100000: color_data = 12'b111111111111;
		12'b011010100001: color_data = 12'b111111111111;
		12'b011010100010: color_data = 12'b111111111111;
		12'b011010100011: color_data = 12'b111111111111;
		12'b011010100100: color_data = 12'b000000000000;
		12'b011010100101: color_data = 12'b111111111111;
		12'b011010100110: color_data = 12'b111111111111;
		12'b011010100111: color_data = 12'b111111111111;
		12'b011010101000: color_data = 12'b111111111111;
		12'b011010101001: color_data = 12'b111111111111;
		12'b011010101010: color_data = 12'b000000000000;
		12'b011010101011: color_data = 12'b111111111111;
		12'b011010101100: color_data = 12'b111111111111;
		12'b011010101101: color_data = 12'b111111111111;
		12'b011010101110: color_data = 12'b111111111111;
		12'b011010101111: color_data = 12'b111111111111;

		12'b011010110000: color_data = 12'b111111111111;
		12'b011010110001: color_data = 12'b111111111111;
		12'b011010110010: color_data = 12'b111111111111;
		12'b011010110011: color_data = 12'b111111111111;
		12'b011010110100: color_data = 12'b000000000000;
		12'b011010110101: color_data = 12'b111111111111;
		12'b011010110110: color_data = 12'b111111111111;
		12'b011010110111: color_data = 12'b111111111111;
		12'b011010111000: color_data = 12'b111111111111;
		12'b011010111001: color_data = 12'b111111111111;
		12'b011010111010: color_data = 12'b000000000000;
		12'b011010111011: color_data = 12'b111111111111;
		12'b011010111100: color_data = 12'b111111111111;
		12'b011010111101: color_data = 12'b111111111111;
		12'b011010111110: color_data = 12'b111111111111;
		12'b011010111111: color_data = 12'b111111111111;

		12'b011011000000: color_data = 12'b111111111111;
		12'b011011000001: color_data = 12'b111111111111;
		12'b011011000010: color_data = 12'b111111111111;
		12'b011011000011: color_data = 12'b111111111111;
		12'b011011000100: color_data = 12'b000000000000;
		12'b011011000101: color_data = 12'b111111111111;
		12'b011011000110: color_data = 12'b111111111111;
		12'b011011000111: color_data = 12'b111111111111;
		12'b011011001000: color_data = 12'b111111111111;
		12'b011011001001: color_data = 12'b111111111111;
		12'b011011001010: color_data = 12'b000000000000;
		12'b011011001011: color_data = 12'b111111111111;
		12'b011011001100: color_data = 12'b111111111111;
		12'b011011001101: color_data = 12'b111111111111;
		12'b011011001110: color_data = 12'b111111111111;
		12'b011011001111: color_data = 12'b111111111111;

		12'b011011010000: color_data = 12'b111111111111;
		12'b011011010001: color_data = 12'b111111111111;
		12'b011011010010: color_data = 12'b111111111111;
		12'b011011010011: color_data = 12'b111111111111;
		12'b011011010100: color_data = 12'b000000000000;
		12'b011011010101: color_data = 12'b000000000000;
		12'b011011010110: color_data = 12'b000000000000;
		12'b011011010111: color_data = 12'b000000000000;
		12'b011011011000: color_data = 12'b000000000000;
		12'b011011011001: color_data = 12'b000000000000;
		12'b011011011010: color_data = 12'b000000000000;
		12'b011011011011: color_data = 12'b111111111111;
		12'b011011011100: color_data = 12'b111111111111;
		12'b011011011101: color_data = 12'b111111111111;
		12'b011011011110: color_data = 12'b111111111111;
		12'b011011011111: color_data = 12'b111111111111;

		12'b011011100000: color_data = 12'b111111111111;
		12'b011011100001: color_data = 12'b111111111111;
		12'b011011100010: color_data = 12'b111111111111;
		12'b011011100011: color_data = 12'b111111111111;
		12'b011011100100: color_data = 12'b111111111111;
		12'b011011100101: color_data = 12'b111111111111;
		12'b011011100110: color_data = 12'b111111111111;
		12'b011011100111: color_data = 12'b111111111111;
		12'b011011101000: color_data = 12'b111111111111;
		12'b011011101001: color_data = 12'b111111111111;
		12'b011011101010: color_data = 12'b111111111111;
		12'b011011101011: color_data = 12'b111111111111;
		12'b011011101100: color_data = 12'b111111111111;
		12'b011011101101: color_data = 12'b111111111111;
		12'b011011101110: color_data = 12'b111111111111;
		12'b011011101111: color_data = 12'b111111111111;

		12'b011011110000: color_data = 12'b111111111111;
		12'b011011110001: color_data = 12'b111111111111;
		12'b011011110010: color_data = 12'b111111111111;
		12'b011011110011: color_data = 12'b111111111111;
		12'b011011110100: color_data = 12'b111111111111;
		12'b011011110101: color_data = 12'b111111111111;
		12'b011011110110: color_data = 12'b111111111111;
		12'b011011110111: color_data = 12'b111111111111;
		12'b011011111000: color_data = 12'b111111111111;
		12'b011011111001: color_data = 12'b111111111111;
		12'b011011111010: color_data = 12'b111111111111;
		12'b011011111011: color_data = 12'b111111111111;
		12'b011011111100: color_data = 12'b111111111111;
		12'b011011111101: color_data = 12'b111111111111;
		12'b011011111110: color_data = 12'b111111111111;
		12'b011011111111: color_data = 12'b111111111111;

		12'b011100000000: color_data = 12'b111111111111;
		12'b011100000001: color_data = 12'b111111111111;
		12'b011100000010: color_data = 12'b111111111111;
		12'b011100000011: color_data = 12'b111111111111;
		12'b011100000100: color_data = 12'b111111111111;
		12'b011100000101: color_data = 12'b111111111111;
		12'b011100000110: color_data = 12'b111111111111;
		12'b011100000111: color_data = 12'b111111111111;
		12'b011100001000: color_data = 12'b111111111111;
		12'b011100001001: color_data = 12'b111111111111;
		12'b011100001010: color_data = 12'b111111111111;
		12'b011100001011: color_data = 12'b111111111111;
		12'b011100001100: color_data = 12'b111111111111;
		12'b011100001101: color_data = 12'b111111111111;
		12'b011100001110: color_data = 12'b111111111111;
		12'b011100001111: color_data = 12'b111111111111;

		12'b011100010000: color_data = 12'b111111111111;
		12'b011100010001: color_data = 12'b111111111111;
		12'b011100010010: color_data = 12'b111111111111;
		12'b011100010011: color_data = 12'b111111111111;
		12'b011100010100: color_data = 12'b000000000000;
		12'b011100010101: color_data = 12'b000000000000;
		12'b011100010110: color_data = 12'b000000000000;
		12'b011100010111: color_data = 12'b000000000000;
		12'b011100011000: color_data = 12'b000000000000;
		12'b011100011001: color_data = 12'b000000000000;
		12'b011100011010: color_data = 12'b000000000000;
		12'b011100011011: color_data = 12'b111111111111;
		12'b011100011100: color_data = 12'b111111111111;
		12'b011100011101: color_data = 12'b111111111111;
		12'b011100011110: color_data = 12'b111111111111;
		12'b011100011111: color_data = 12'b111111111111;

		12'b011100100000: color_data = 12'b111111111111;
		12'b011100100001: color_data = 12'b111111111111;
		12'b011100100010: color_data = 12'b111111111111;
		12'b011100100011: color_data = 12'b111111111111;
		12'b011100100100: color_data = 12'b000000000000;
		12'b011100100101: color_data = 12'b111111111111;
		12'b011100100110: color_data = 12'b111111111111;
		12'b011100100111: color_data = 12'b111111111111;
		12'b011100101000: color_data = 12'b111111111111;
		12'b011100101001: color_data = 12'b111111111111;
		12'b011100101010: color_data = 12'b000000000000;
		12'b011100101011: color_data = 12'b111111111111;
		12'b011100101100: color_data = 12'b111111111111;
		12'b011100101101: color_data = 12'b111111111111;
		12'b011100101110: color_data = 12'b111111111111;
		12'b011100101111: color_data = 12'b111111111111;

		12'b011100110000: color_data = 12'b111111111111;
		12'b011100110001: color_data = 12'b111111111111;
		12'b011100110010: color_data = 12'b111111111111;
		12'b011100110011: color_data = 12'b111111111111;
		12'b011100110100: color_data = 12'b000000000000;
		12'b011100110101: color_data = 12'b111111111111;
		12'b011100110110: color_data = 12'b111111111111;
		12'b011100110111: color_data = 12'b111111111111;
		12'b011100111000: color_data = 12'b111111111111;
		12'b011100111001: color_data = 12'b111111111111;
		12'b011100111010: color_data = 12'b000000000000;
		12'b011100111011: color_data = 12'b111111111111;
		12'b011100111100: color_data = 12'b111111111111;
		12'b011100111101: color_data = 12'b111111111111;
		12'b011100111110: color_data = 12'b111111111111;
		12'b011100111111: color_data = 12'b111111111111;

		12'b011101000000: color_data = 12'b111111111111;
		12'b011101000001: color_data = 12'b111111111111;
		12'b011101000010: color_data = 12'b111111111111;
		12'b011101000011: color_data = 12'b111111111111;
		12'b011101000100: color_data = 12'b111111111111;
		12'b011101000101: color_data = 12'b111111111111;
		12'b011101000110: color_data = 12'b111111111111;
		12'b011101000111: color_data = 12'b111111111111;
		12'b011101001000: color_data = 12'b111111111111;
		12'b011101001001: color_data = 12'b111111111111;
		12'b011101001010: color_data = 12'b000000000000;
		12'b011101001011: color_data = 12'b111111111111;
		12'b011101001100: color_data = 12'b111111111111;
		12'b011101001101: color_data = 12'b111111111111;
		12'b011101001110: color_data = 12'b111111111111;
		12'b011101001111: color_data = 12'b111111111111;

		12'b011101010000: color_data = 12'b111111111111;
		12'b011101010001: color_data = 12'b111111111111;
		12'b011101010010: color_data = 12'b111111111111;
		12'b011101010011: color_data = 12'b111111111111;
		12'b011101010100: color_data = 12'b111111111111;
		12'b011101010101: color_data = 12'b111111111111;
		12'b011101010110: color_data = 12'b111111111111;
		12'b011101010111: color_data = 12'b111111111111;
		12'b011101011000: color_data = 12'b111111111111;
		12'b011101011001: color_data = 12'b111111111111;
		12'b011101011010: color_data = 12'b000000000000;
		12'b011101011011: color_data = 12'b111111111111;
		12'b011101011100: color_data = 12'b111111111111;
		12'b011101011101: color_data = 12'b111111111111;
		12'b011101011110: color_data = 12'b111111111111;
		12'b011101011111: color_data = 12'b111111111111;

		12'b011101100000: color_data = 12'b111111111111;
		12'b011101100001: color_data = 12'b111111111111;
		12'b011101100010: color_data = 12'b111111111111;
		12'b011101100011: color_data = 12'b111111111111;
		12'b011101100100: color_data = 12'b111111111111;
		12'b011101100101: color_data = 12'b111111111111;
		12'b011101100110: color_data = 12'b111111111111;
		12'b011101100111: color_data = 12'b111111111111;
		12'b011101101000: color_data = 12'b111111111111;
		12'b011101101001: color_data = 12'b111111111111;
		12'b011101101010: color_data = 12'b000000000000;
		12'b011101101011: color_data = 12'b111111111111;
		12'b011101101100: color_data = 12'b111111111111;
		12'b011101101101: color_data = 12'b111111111111;
		12'b011101101110: color_data = 12'b111111111111;
		12'b011101101111: color_data = 12'b111111111111;

		12'b011101110000: color_data = 12'b111111111111;
		12'b011101110001: color_data = 12'b111111111111;
		12'b011101110010: color_data = 12'b111111111111;
		12'b011101110011: color_data = 12'b111111111111;
		12'b011101110100: color_data = 12'b111111111111;
		12'b011101110101: color_data = 12'b111111111111;
		12'b011101110110: color_data = 12'b111111111111;
		12'b011101110111: color_data = 12'b111111111111;
		12'b011101111000: color_data = 12'b000000000000;
		12'b011101111001: color_data = 12'b000000000000;
		12'b011101111010: color_data = 12'b000000000000;
		12'b011101111011: color_data = 12'b111111111111;
		12'b011101111100: color_data = 12'b111111111111;
		12'b011101111101: color_data = 12'b111111111111;
		12'b011101111110: color_data = 12'b111111111111;
		12'b011101111111: color_data = 12'b111111111111;

		12'b011110000000: color_data = 12'b111111111111;
		12'b011110000001: color_data = 12'b111111111111;
		12'b011110000010: color_data = 12'b111111111111;
		12'b011110000011: color_data = 12'b111111111111;
		12'b011110000100: color_data = 12'b111111111111;
		12'b011110000101: color_data = 12'b111111111111;
		12'b011110000110: color_data = 12'b111111111111;
		12'b011110000111: color_data = 12'b111111111111;
		12'b011110001000: color_data = 12'b000000000000;
		12'b011110001001: color_data = 12'b111111111111;
		12'b011110001010: color_data = 12'b111111111111;
		12'b011110001011: color_data = 12'b111111111111;
		12'b011110001100: color_data = 12'b111111111111;
		12'b011110001101: color_data = 12'b111111111111;
		12'b011110001110: color_data = 12'b111111111111;
		12'b011110001111: color_data = 12'b111111111111;

		12'b011110010000: color_data = 12'b111111111111;
		12'b011110010001: color_data = 12'b111111111111;
		12'b011110010010: color_data = 12'b111111111111;
		12'b011110010011: color_data = 12'b111111111111;
		12'b011110010100: color_data = 12'b111111111111;
		12'b011110010101: color_data = 12'b111111111111;
		12'b011110010110: color_data = 12'b111111111111;
		12'b011110010111: color_data = 12'b111111111111;
		12'b011110011000: color_data = 12'b000000000000;
		12'b011110011001: color_data = 12'b111111111111;
		12'b011110011010: color_data = 12'b111111111111;
		12'b011110011011: color_data = 12'b111111111111;
		12'b011110011100: color_data = 12'b111111111111;
		12'b011110011101: color_data = 12'b111111111111;
		12'b011110011110: color_data = 12'b111111111111;
		12'b011110011111: color_data = 12'b111111111111;

		12'b011110100000: color_data = 12'b111111111111;
		12'b011110100001: color_data = 12'b111111111111;
		12'b011110100010: color_data = 12'b111111111111;
		12'b011110100011: color_data = 12'b111111111111;
		12'b011110100100: color_data = 12'b111111111111;
		12'b011110100101: color_data = 12'b111111111111;
		12'b011110100110: color_data = 12'b111111111111;
		12'b011110100111: color_data = 12'b111111111111;
		12'b011110101000: color_data = 12'b000000000000;
		12'b011110101001: color_data = 12'b111111111111;
		12'b011110101010: color_data = 12'b111111111111;
		12'b011110101011: color_data = 12'b111111111111;
		12'b011110101100: color_data = 12'b111111111111;
		12'b011110101101: color_data = 12'b111111111111;
		12'b011110101110: color_data = 12'b111111111111;
		12'b011110101111: color_data = 12'b111111111111;

		12'b011110110000: color_data = 12'b111111111111;
		12'b011110110001: color_data = 12'b111111111111;
		12'b011110110010: color_data = 12'b111111111111;
		12'b011110110011: color_data = 12'b111111111111;
		12'b011110110100: color_data = 12'b111111111111;
		12'b011110110101: color_data = 12'b111111111111;
		12'b011110110110: color_data = 12'b111111111111;
		12'b011110110111: color_data = 12'b111111111111;
		12'b011110111000: color_data = 12'b000000000000;
		12'b011110111001: color_data = 12'b111111111111;
		12'b011110111010: color_data = 12'b111111111111;
		12'b011110111011: color_data = 12'b111111111111;
		12'b011110111100: color_data = 12'b111111111111;
		12'b011110111101: color_data = 12'b111111111111;
		12'b011110111110: color_data = 12'b111111111111;
		12'b011110111111: color_data = 12'b111111111111;

		12'b011111000000: color_data = 12'b111111111111;
		12'b011111000001: color_data = 12'b111111111111;
		12'b011111000010: color_data = 12'b111111111111;
		12'b011111000011: color_data = 12'b111111111111;
		12'b011111000100: color_data = 12'b111111111111;
		12'b011111000101: color_data = 12'b111111111111;
		12'b011111000110: color_data = 12'b111111111111;
		12'b011111000111: color_data = 12'b111111111111;
		12'b011111001000: color_data = 12'b000000000000;
		12'b011111001001: color_data = 12'b111111111111;
		12'b011111001010: color_data = 12'b111111111111;
		12'b011111001011: color_data = 12'b111111111111;
		12'b011111001100: color_data = 12'b111111111111;
		12'b011111001101: color_data = 12'b111111111111;
		12'b011111001110: color_data = 12'b111111111111;
		12'b011111001111: color_data = 12'b111111111111;

		12'b011111010000: color_data = 12'b111111111111;
		12'b011111010001: color_data = 12'b111111111111;
		12'b011111010010: color_data = 12'b111111111111;
		12'b011111010011: color_data = 12'b111111111111;
		12'b011111010100: color_data = 12'b111111111111;
		12'b011111010101: color_data = 12'b111111111111;
		12'b011111010110: color_data = 12'b111111111111;
		12'b011111010111: color_data = 12'b111111111111;
		12'b011111011000: color_data = 12'b000000000000;
		12'b011111011001: color_data = 12'b111111111111;
		12'b011111011010: color_data = 12'b111111111111;
		12'b011111011011: color_data = 12'b111111111111;
		12'b011111011100: color_data = 12'b111111111111;
		12'b011111011101: color_data = 12'b111111111111;
		12'b011111011110: color_data = 12'b111111111111;
		12'b011111011111: color_data = 12'b111111111111;

		12'b011111100000: color_data = 12'b111111111111;
		12'b011111100001: color_data = 12'b111111111111;
		12'b011111100010: color_data = 12'b111111111111;
		12'b011111100011: color_data = 12'b111111111111;
		12'b011111100100: color_data = 12'b111111111111;
		12'b011111100101: color_data = 12'b111111111111;
		12'b011111100110: color_data = 12'b111111111111;
		12'b011111100111: color_data = 12'b111111111111;
		12'b011111101000: color_data = 12'b111111111111;
		12'b011111101001: color_data = 12'b111111111111;
		12'b011111101010: color_data = 12'b111111111111;
		12'b011111101011: color_data = 12'b111111111111;
		12'b011111101100: color_data = 12'b111111111111;
		12'b011111101101: color_data = 12'b111111111111;
		12'b011111101110: color_data = 12'b111111111111;
		12'b011111101111: color_data = 12'b111111111111;

		12'b011111110000: color_data = 12'b111111111111;
		12'b011111110001: color_data = 12'b111111111111;
		12'b011111110010: color_data = 12'b111111111111;
		12'b011111110011: color_data = 12'b111111111111;
		12'b011111110100: color_data = 12'b111111111111;
		12'b011111110101: color_data = 12'b111111111111;
		12'b011111110110: color_data = 12'b111111111111;
		12'b011111110111: color_data = 12'b111111111111;
		12'b011111111000: color_data = 12'b111111111111;
		12'b011111111001: color_data = 12'b111111111111;
		12'b011111111010: color_data = 12'b111111111111;
		12'b011111111011: color_data = 12'b111111111111;
		12'b011111111100: color_data = 12'b111111111111;
		12'b011111111101: color_data = 12'b111111111111;
		12'b011111111110: color_data = 12'b111111111111;
		12'b011111111111: color_data = 12'b111111111111;

		12'b100000000000: color_data = 12'b111111111111;
		12'b100000000001: color_data = 12'b111111111111;
		12'b100000000010: color_data = 12'b111111111111;
		12'b100000000011: color_data = 12'b111111111111;
		12'b100000000100: color_data = 12'b111111111111;
		12'b100000000101: color_data = 12'b111111111111;
		12'b100000000110: color_data = 12'b111111111111;
		12'b100000000111: color_data = 12'b111111111111;
		12'b100000001000: color_data = 12'b111111111111;
		12'b100000001001: color_data = 12'b111111111111;
		12'b100000001010: color_data = 12'b111111111111;
		12'b100000001011: color_data = 12'b111111111111;
		12'b100000001100: color_data = 12'b111111111111;
		12'b100000001101: color_data = 12'b111111111111;
		12'b100000001110: color_data = 12'b111111111111;
		12'b100000001111: color_data = 12'b111111111111;

		12'b100000010000: color_data = 12'b111111111111;
		12'b100000010001: color_data = 12'b111111111111;
		12'b100000010010: color_data = 12'b111111111111;
		12'b100000010011: color_data = 12'b111111111111;
		12'b100000010100: color_data = 12'b000000000000;
		12'b100000010101: color_data = 12'b000000000000;
		12'b100000010110: color_data = 12'b000000000000;
		12'b100000010111: color_data = 12'b000000000000;
		12'b100000011000: color_data = 12'b000000000000;
		12'b100000011001: color_data = 12'b000000000000;
		12'b100000011010: color_data = 12'b000000000000;
		12'b100000011011: color_data = 12'b111111111111;
		12'b100000011100: color_data = 12'b111111111111;
		12'b100000011101: color_data = 12'b111111111111;
		12'b100000011110: color_data = 12'b111111111111;
		12'b100000011111: color_data = 12'b111111111111;

		12'b100000100000: color_data = 12'b111111111111;
		12'b100000100001: color_data = 12'b111111111111;
		12'b100000100010: color_data = 12'b111111111111;
		12'b100000100011: color_data = 12'b111111111111;
		12'b100000100100: color_data = 12'b000000000000;
		12'b100000100101: color_data = 12'b111111111111;
		12'b100000100110: color_data = 12'b111111111111;
		12'b100000100111: color_data = 12'b111111111111;
		12'b100000101000: color_data = 12'b111111111111;
		12'b100000101001: color_data = 12'b111111111111;
		12'b100000101010: color_data = 12'b000000000000;
		12'b100000101011: color_data = 12'b111111111111;
		12'b100000101100: color_data = 12'b111111111111;
		12'b100000101101: color_data = 12'b111111111111;
		12'b100000101110: color_data = 12'b111111111111;
		12'b100000101111: color_data = 12'b111111111111;

		12'b100000110000: color_data = 12'b111111111111;
		12'b100000110001: color_data = 12'b111111111111;
		12'b100000110010: color_data = 12'b111111111111;
		12'b100000110011: color_data = 12'b111111111111;
		12'b100000110100: color_data = 12'b000000000000;
		12'b100000110101: color_data = 12'b111111111111;
		12'b100000110110: color_data = 12'b111111111111;
		12'b100000110111: color_data = 12'b111111111111;
		12'b100000111000: color_data = 12'b111111111111;
		12'b100000111001: color_data = 12'b111111111111;
		12'b100000111010: color_data = 12'b000000000000;
		12'b100000111011: color_data = 12'b111111111111;
		12'b100000111100: color_data = 12'b111111111111;
		12'b100000111101: color_data = 12'b111111111111;
		12'b100000111110: color_data = 12'b111111111111;
		12'b100000111111: color_data = 12'b111111111111;

		12'b100001000000: color_data = 12'b111111111111;
		12'b100001000001: color_data = 12'b111111111111;
		12'b100001000010: color_data = 12'b111111111111;
		12'b100001000011: color_data = 12'b111111111111;
		12'b100001000100: color_data = 12'b000000000000;
		12'b100001000101: color_data = 12'b111111111111;
		12'b100001000110: color_data = 12'b111111111111;
		12'b100001000111: color_data = 12'b111111111111;
		12'b100001001000: color_data = 12'b111111111111;
		12'b100001001001: color_data = 12'b111111111111;
		12'b100001001010: color_data = 12'b000000000000;
		12'b100001001011: color_data = 12'b111111111111;
		12'b100001001100: color_data = 12'b111111111111;
		12'b100001001101: color_data = 12'b111111111111;
		12'b100001001110: color_data = 12'b111111111111;
		12'b100001001111: color_data = 12'b111111111111;

		12'b100001010000: color_data = 12'b111111111111;
		12'b100001010001: color_data = 12'b111111111111;
		12'b100001010010: color_data = 12'b111111111111;
		12'b100001010011: color_data = 12'b111111111111;
		12'b100001010100: color_data = 12'b000000000000;
		12'b100001010101: color_data = 12'b111111111111;
		12'b100001010110: color_data = 12'b111111111111;
		12'b100001010111: color_data = 12'b111111111111;
		12'b100001011000: color_data = 12'b111111111111;
		12'b100001011001: color_data = 12'b111111111111;
		12'b100001011010: color_data = 12'b000000000000;
		12'b100001011011: color_data = 12'b111111111111;
		12'b100001011100: color_data = 12'b111111111111;
		12'b100001011101: color_data = 12'b111111111111;
		12'b100001011110: color_data = 12'b111111111111;
		12'b100001011111: color_data = 12'b111111111111;

		12'b100001100000: color_data = 12'b111111111111;
		12'b100001100001: color_data = 12'b111111111111;
		12'b100001100010: color_data = 12'b111111111111;
		12'b100001100011: color_data = 12'b111111111111;
		12'b100001100100: color_data = 12'b000000000000;
		12'b100001100101: color_data = 12'b111111111111;
		12'b100001100110: color_data = 12'b111111111111;
		12'b100001100111: color_data = 12'b111111111111;
		12'b100001101000: color_data = 12'b111111111111;
		12'b100001101001: color_data = 12'b111111111111;
		12'b100001101010: color_data = 12'b000000000000;
		12'b100001101011: color_data = 12'b111111111111;
		12'b100001101100: color_data = 12'b111111111111;
		12'b100001101101: color_data = 12'b111111111111;
		12'b100001101110: color_data = 12'b111111111111;
		12'b100001101111: color_data = 12'b111111111111;

		12'b100001110000: color_data = 12'b111111111111;
		12'b100001110001: color_data = 12'b111111111111;
		12'b100001110010: color_data = 12'b111111111111;
		12'b100001110011: color_data = 12'b111111111111;
		12'b100001110100: color_data = 12'b000000000000;
		12'b100001110101: color_data = 12'b111111111111;
		12'b100001110110: color_data = 12'b111111111111;
		12'b100001110111: color_data = 12'b111111111111;
		12'b100001111000: color_data = 12'b111111111111;
		12'b100001111001: color_data = 12'b111111111111;
		12'b100001111010: color_data = 12'b000000000000;
		12'b100001111011: color_data = 12'b111111111111;
		12'b100001111100: color_data = 12'b111111111111;
		12'b100001111101: color_data = 12'b111111111111;
		12'b100001111110: color_data = 12'b111111111111;
		12'b100001111111: color_data = 12'b111111111111;

		12'b100010000000: color_data = 12'b111111111111;
		12'b100010000001: color_data = 12'b111111111111;
		12'b100010000010: color_data = 12'b111111111111;
		12'b100010000011: color_data = 12'b111111111111;
		12'b100010000100: color_data = 12'b000000000000;
		12'b100010000101: color_data = 12'b000000000000;
		12'b100010000110: color_data = 12'b000000000000;
		12'b100010000111: color_data = 12'b000000000000;
		12'b100010001000: color_data = 12'b000000000000;
		12'b100010001001: color_data = 12'b000000000000;
		12'b100010001010: color_data = 12'b000000000000;
		12'b100010001011: color_data = 12'b111111111111;
		12'b100010001100: color_data = 12'b111111111111;
		12'b100010001101: color_data = 12'b111111111111;
		12'b100010001110: color_data = 12'b111111111111;
		12'b100010001111: color_data = 12'b111111111111;

		12'b100010010000: color_data = 12'b111111111111;
		12'b100010010001: color_data = 12'b111111111111;
		12'b100010010010: color_data = 12'b111111111111;
		12'b100010010011: color_data = 12'b111111111111;
		12'b100010010100: color_data = 12'b000000000000;
		12'b100010010101: color_data = 12'b111111111111;
		12'b100010010110: color_data = 12'b111111111111;
		12'b100010010111: color_data = 12'b111111111111;
		12'b100010011000: color_data = 12'b111111111111;
		12'b100010011001: color_data = 12'b111111111111;
		12'b100010011010: color_data = 12'b000000000000;
		12'b100010011011: color_data = 12'b111111111111;
		12'b100010011100: color_data = 12'b111111111111;
		12'b100010011101: color_data = 12'b111111111111;
		12'b100010011110: color_data = 12'b111111111111;
		12'b100010011111: color_data = 12'b111111111111;

		12'b100010100000: color_data = 12'b111111111111;
		12'b100010100001: color_data = 12'b111111111111;
		12'b100010100010: color_data = 12'b111111111111;
		12'b100010100011: color_data = 12'b111111111111;
		12'b100010100100: color_data = 12'b000000000000;
		12'b100010100101: color_data = 12'b111111111111;
		12'b100010100110: color_data = 12'b111111111111;
		12'b100010100111: color_data = 12'b111111111111;
		12'b100010101000: color_data = 12'b111111111111;
		12'b100010101001: color_data = 12'b111111111111;
		12'b100010101010: color_data = 12'b000000000000;
		12'b100010101011: color_data = 12'b111111111111;
		12'b100010101100: color_data = 12'b111111111111;
		12'b100010101101: color_data = 12'b111111111111;
		12'b100010101110: color_data = 12'b111111111111;
		12'b100010101111: color_data = 12'b111111111111;

		12'b100010110000: color_data = 12'b111111111111;
		12'b100010110001: color_data = 12'b111111111111;
		12'b100010110010: color_data = 12'b111111111111;
		12'b100010110011: color_data = 12'b111111111111;
		12'b100010110100: color_data = 12'b000000000000;
		12'b100010110101: color_data = 12'b111111111111;
		12'b100010110110: color_data = 12'b111111111111;
		12'b100010110111: color_data = 12'b111111111111;
		12'b100010111000: color_data = 12'b111111111111;
		12'b100010111001: color_data = 12'b111111111111;
		12'b100010111010: color_data = 12'b000000000000;
		12'b100010111011: color_data = 12'b111111111111;
		12'b100010111100: color_data = 12'b111111111111;
		12'b100010111101: color_data = 12'b111111111111;
		12'b100010111110: color_data = 12'b111111111111;
		12'b100010111111: color_data = 12'b111111111111;

		12'b100011000000: color_data = 12'b111111111111;
		12'b100011000001: color_data = 12'b111111111111;
		12'b100011000010: color_data = 12'b111111111111;
		12'b100011000011: color_data = 12'b111111111111;
		12'b100011000100: color_data = 12'b000000000000;
		12'b100011000101: color_data = 12'b111111111111;
		12'b100011000110: color_data = 12'b111111111111;
		12'b100011000111: color_data = 12'b111111111111;
		12'b100011001000: color_data = 12'b111111111111;
		12'b100011001001: color_data = 12'b111111111111;
		12'b100011001010: color_data = 12'b000000000000;
		12'b100011001011: color_data = 12'b111111111111;
		12'b100011001100: color_data = 12'b111111111111;
		12'b100011001101: color_data = 12'b111111111111;
		12'b100011001110: color_data = 12'b111111111111;
		12'b100011001111: color_data = 12'b111111111111;

		12'b100011010000: color_data = 12'b111111111111;
		12'b100011010001: color_data = 12'b111111111111;
		12'b100011010010: color_data = 12'b111111111111;
		12'b100011010011: color_data = 12'b111111111111;
		12'b100011010100: color_data = 12'b000000000000;
		12'b100011010101: color_data = 12'b000000000000;
		12'b100011010110: color_data = 12'b000000000000;
		12'b100011010111: color_data = 12'b000000000000;
		12'b100011011000: color_data = 12'b000000000000;
		12'b100011011001: color_data = 12'b000000000000;
		12'b100011011010: color_data = 12'b000000000000;
		12'b100011011011: color_data = 12'b111111111111;
		12'b100011011100: color_data = 12'b111111111111;
		12'b100011011101: color_data = 12'b111111111111;
		12'b100011011110: color_data = 12'b111111111111;
		12'b100011011111: color_data = 12'b111111111111;

		12'b100011100000: color_data = 12'b111111111111;
		12'b100011100001: color_data = 12'b111111111111;
		12'b100011100010: color_data = 12'b111111111111;
		12'b100011100011: color_data = 12'b111111111111;
		12'b100011100100: color_data = 12'b111111111111;
		12'b100011100101: color_data = 12'b111111111111;
		12'b100011100110: color_data = 12'b111111111111;
		12'b100011100111: color_data = 12'b111111111111;
		12'b100011101000: color_data = 12'b111111111111;
		12'b100011101001: color_data = 12'b111111111111;
		12'b100011101010: color_data = 12'b111111111111;
		12'b100011101011: color_data = 12'b111111111111;
		12'b100011101100: color_data = 12'b111111111111;
		12'b100011101101: color_data = 12'b111111111111;
		12'b100011101110: color_data = 12'b111111111111;
		12'b100011101111: color_data = 12'b111111111111;

		12'b100011110000: color_data = 12'b111111111111;
		12'b100011110001: color_data = 12'b111111111111;
		12'b100011110010: color_data = 12'b111111111111;
		12'b100011110011: color_data = 12'b111111111111;
		12'b100011110100: color_data = 12'b111111111111;
		12'b100011110101: color_data = 12'b111111111111;
		12'b100011110110: color_data = 12'b111111111111;
		12'b100011110111: color_data = 12'b111111111111;
		12'b100011111000: color_data = 12'b111111111111;
		12'b100011111001: color_data = 12'b111111111111;
		12'b100011111010: color_data = 12'b111111111111;
		12'b100011111011: color_data = 12'b111111111111;
		12'b100011111100: color_data = 12'b111111111111;
		12'b100011111101: color_data = 12'b111111111111;
		12'b100011111110: color_data = 12'b111111111111;
		12'b100011111111: color_data = 12'b111111111111;

		12'b100100000000: color_data = 12'b111111111111;
		12'b100100000001: color_data = 12'b111111111111;
		12'b100100000010: color_data = 12'b111111111111;
		12'b100100000011: color_data = 12'b111111111111;
		12'b100100000100: color_data = 12'b111111111111;
		12'b100100000101: color_data = 12'b111111111111;
		12'b100100000110: color_data = 12'b111111111111;
		12'b100100000111: color_data = 12'b111111111111;
		12'b100100001000: color_data = 12'b111111111111;
		12'b100100001001: color_data = 12'b111111111111;
		12'b100100001010: color_data = 12'b111111111111;
		12'b100100001011: color_data = 12'b111111111111;
		12'b100100001100: color_data = 12'b111111111111;
		12'b100100001101: color_data = 12'b111111111111;
		12'b100100001110: color_data = 12'b111111111111;
		12'b100100001111: color_data = 12'b111111111111;

		12'b100100010000: color_data = 12'b111111111111;
		12'b100100010001: color_data = 12'b111111111111;
		12'b100100010010: color_data = 12'b111111111111;
		12'b100100010011: color_data = 12'b111111111111;
		12'b100100010100: color_data = 12'b000000000000;
		12'b100100010101: color_data = 12'b000000000000;
		12'b100100010110: color_data = 12'b000000000000;
		12'b100100010111: color_data = 12'b000000000000;
		12'b100100011000: color_data = 12'b000000000000;
		12'b100100011001: color_data = 12'b000000000000;
		12'b100100011010: color_data = 12'b000000000000;
		12'b100100011011: color_data = 12'b111111111111;
		12'b100100011100: color_data = 12'b111111111111;
		12'b100100011101: color_data = 12'b111111111111;
		12'b100100011110: color_data = 12'b111111111111;
		12'b100100011111: color_data = 12'b111111111111;

		12'b100100100000: color_data = 12'b111111111111;
		12'b100100100001: color_data = 12'b111111111111;
		12'b100100100010: color_data = 12'b111111111111;
		12'b100100100011: color_data = 12'b111111111111;
		12'b100100100100: color_data = 12'b000000000000;
		12'b100100100101: color_data = 12'b111111111111;
		12'b100100100110: color_data = 12'b111111111111;
		12'b100100100111: color_data = 12'b111111111111;
		12'b100100101000: color_data = 12'b111111111111;
		12'b100100101001: color_data = 12'b111111111111;
		12'b100100101010: color_data = 12'b000000000000;
		12'b100100101011: color_data = 12'b111111111111;
		12'b100100101100: color_data = 12'b111111111111;
		12'b100100101101: color_data = 12'b111111111111;
		12'b100100101110: color_data = 12'b111111111111;
		12'b100100101111: color_data = 12'b111111111111;

		12'b100100110000: color_data = 12'b111111111111;
		12'b100100110001: color_data = 12'b111111111111;
		12'b100100110010: color_data = 12'b111111111111;
		12'b100100110011: color_data = 12'b111111111111;
		12'b100100110100: color_data = 12'b000000000000;
		12'b100100110101: color_data = 12'b111111111111;
		12'b100100110110: color_data = 12'b111111111111;
		12'b100100110111: color_data = 12'b111111111111;
		12'b100100111000: color_data = 12'b111111111111;
		12'b100100111001: color_data = 12'b111111111111;
		12'b100100111010: color_data = 12'b000000000000;
		12'b100100111011: color_data = 12'b111111111111;
		12'b100100111100: color_data = 12'b111111111111;
		12'b100100111101: color_data = 12'b111111111111;
		12'b100100111110: color_data = 12'b111111111111;
		12'b100100111111: color_data = 12'b111111111111;

		12'b100101000000: color_data = 12'b111111111111;
		12'b100101000001: color_data = 12'b111111111111;
		12'b100101000010: color_data = 12'b111111111111;
		12'b100101000011: color_data = 12'b111111111111;
		12'b100101000100: color_data = 12'b000000000000;
		12'b100101000101: color_data = 12'b111111111111;
		12'b100101000110: color_data = 12'b111111111111;
		12'b100101000111: color_data = 12'b111111111111;
		12'b100101001000: color_data = 12'b111111111111;
		12'b100101001001: color_data = 12'b111111111111;
		12'b100101001010: color_data = 12'b000000000000;
		12'b100101001011: color_data = 12'b111111111111;
		12'b100101001100: color_data = 12'b111111111111;
		12'b100101001101: color_data = 12'b111111111111;
		12'b100101001110: color_data = 12'b111111111111;
		12'b100101001111: color_data = 12'b111111111111;

		12'b100101010000: color_data = 12'b111111111111;
		12'b100101010001: color_data = 12'b111111111111;
		12'b100101010010: color_data = 12'b111111111111;
		12'b100101010011: color_data = 12'b111111111111;
		12'b100101010100: color_data = 12'b000000000000;
		12'b100101010101: color_data = 12'b111111111111;
		12'b100101010110: color_data = 12'b111111111111;
		12'b100101010111: color_data = 12'b111111111111;
		12'b100101011000: color_data = 12'b111111111111;
		12'b100101011001: color_data = 12'b111111111111;
		12'b100101011010: color_data = 12'b000000000000;
		12'b100101011011: color_data = 12'b111111111111;
		12'b100101011100: color_data = 12'b111111111111;
		12'b100101011101: color_data = 12'b111111111111;
		12'b100101011110: color_data = 12'b111111111111;
		12'b100101011111: color_data = 12'b111111111111;

		12'b100101100000: color_data = 12'b111111111111;
		12'b100101100001: color_data = 12'b111111111111;
		12'b100101100010: color_data = 12'b111111111111;
		12'b100101100011: color_data = 12'b111111111111;
		12'b100101100100: color_data = 12'b000000000000;
		12'b100101100101: color_data = 12'b111111111111;
		12'b100101100110: color_data = 12'b111111111111;
		12'b100101100111: color_data = 12'b111111111111;
		12'b100101101000: color_data = 12'b111111111111;
		12'b100101101001: color_data = 12'b111111111111;
		12'b100101101010: color_data = 12'b000000000000;
		12'b100101101011: color_data = 12'b111111111111;
		12'b100101101100: color_data = 12'b111111111111;
		12'b100101101101: color_data = 12'b111111111111;
		12'b100101101110: color_data = 12'b111111111111;
		12'b100101101111: color_data = 12'b111111111111;

		12'b100101110000: color_data = 12'b111111111111;
		12'b100101110001: color_data = 12'b111111111111;
		12'b100101110010: color_data = 12'b111111111111;
		12'b100101110011: color_data = 12'b111111111111;
		12'b100101110100: color_data = 12'b000000000000;
		12'b100101110101: color_data = 12'b000000000000;
		12'b100101110110: color_data = 12'b000000000000;
		12'b100101110111: color_data = 12'b000000000000;
		12'b100101111000: color_data = 12'b000000000000;
		12'b100101111001: color_data = 12'b000000000000;
		12'b100101111010: color_data = 12'b000000000000;
		12'b100101111011: color_data = 12'b111111111111;
		12'b100101111100: color_data = 12'b111111111111;
		12'b100101111101: color_data = 12'b111111111111;
		12'b100101111110: color_data = 12'b111111111111;
		12'b100101111111: color_data = 12'b111111111111;

		12'b100110000000: color_data = 12'b111111111111;
		12'b100110000001: color_data = 12'b111111111111;
		12'b100110000010: color_data = 12'b111111111111;
		12'b100110000011: color_data = 12'b111111111111;
		12'b100110000100: color_data = 12'b111111111111;
		12'b100110000101: color_data = 12'b111111111111;
		12'b100110000110: color_data = 12'b111111111111;
		12'b100110000111: color_data = 12'b111111111111;
		12'b100110001000: color_data = 12'b111111111111;
		12'b100110001001: color_data = 12'b111111111111;
		12'b100110001010: color_data = 12'b000000000000;
		12'b100110001011: color_data = 12'b111111111111;
		12'b100110001100: color_data = 12'b111111111111;
		12'b100110001101: color_data = 12'b111111111111;
		12'b100110001110: color_data = 12'b111111111111;
		12'b100110001111: color_data = 12'b111111111111;

		12'b100110010000: color_data = 12'b111111111111;
		12'b100110010001: color_data = 12'b111111111111;
		12'b100110010010: color_data = 12'b111111111111;
		12'b100110010011: color_data = 12'b111111111111;
		12'b100110010100: color_data = 12'b111111111111;
		12'b100110010101: color_data = 12'b111111111111;
		12'b100110010110: color_data = 12'b111111111111;
		12'b100110010111: color_data = 12'b111111111111;
		12'b100110011000: color_data = 12'b111111111111;
		12'b100110011001: color_data = 12'b111111111111;
		12'b100110011010: color_data = 12'b000000000000;
		12'b100110011011: color_data = 12'b111111111111;
		12'b100110011100: color_data = 12'b111111111111;
		12'b100110011101: color_data = 12'b111111111111;
		12'b100110011110: color_data = 12'b111111111111;
		12'b100110011111: color_data = 12'b111111111111;

		12'b100110100000: color_data = 12'b111111111111;
		12'b100110100001: color_data = 12'b111111111111;
		12'b100110100010: color_data = 12'b111111111111;
		12'b100110100011: color_data = 12'b111111111111;
		12'b100110100100: color_data = 12'b111111111111;
		12'b100110100101: color_data = 12'b111111111111;
		12'b100110100110: color_data = 12'b111111111111;
		12'b100110100111: color_data = 12'b111111111111;
		12'b100110101000: color_data = 12'b111111111111;
		12'b100110101001: color_data = 12'b111111111111;
		12'b100110101010: color_data = 12'b000000000000;
		12'b100110101011: color_data = 12'b111111111111;
		12'b100110101100: color_data = 12'b111111111111;
		12'b100110101101: color_data = 12'b111111111111;
		12'b100110101110: color_data = 12'b111111111111;
		12'b100110101111: color_data = 12'b111111111111;

		12'b100110110000: color_data = 12'b111111111111;
		12'b100110110001: color_data = 12'b111111111111;
		12'b100110110010: color_data = 12'b111111111111;
		12'b100110110011: color_data = 12'b111111111111;
		12'b100110110100: color_data = 12'b111111111111;
		12'b100110110101: color_data = 12'b111111111111;
		12'b100110110110: color_data = 12'b111111111111;
		12'b100110110111: color_data = 12'b111111111111;
		12'b100110111000: color_data = 12'b111111111111;
		12'b100110111001: color_data = 12'b111111111111;
		12'b100110111010: color_data = 12'b000000000000;
		12'b100110111011: color_data = 12'b111111111111;
		12'b100110111100: color_data = 12'b111111111111;
		12'b100110111101: color_data = 12'b111111111111;
		12'b100110111110: color_data = 12'b111111111111;
		12'b100110111111: color_data = 12'b111111111111;

		12'b100111000000: color_data = 12'b111111111111;
		12'b100111000001: color_data = 12'b111111111111;
		12'b100111000010: color_data = 12'b111111111111;
		12'b100111000011: color_data = 12'b111111111111;
		12'b100111000100: color_data = 12'b111111111111;
		12'b100111000101: color_data = 12'b111111111111;
		12'b100111000110: color_data = 12'b111111111111;
		12'b100111000111: color_data = 12'b111111111111;
		12'b100111001000: color_data = 12'b111111111111;
		12'b100111001001: color_data = 12'b111111111111;
		12'b100111001010: color_data = 12'b000000000000;
		12'b100111001011: color_data = 12'b111111111111;
		12'b100111001100: color_data = 12'b111111111111;
		12'b100111001101: color_data = 12'b111111111111;
		12'b100111001110: color_data = 12'b111111111111;
		12'b100111001111: color_data = 12'b111111111111;

		12'b100111010000: color_data = 12'b111111111111;
		12'b100111010001: color_data = 12'b111111111111;
		12'b100111010010: color_data = 12'b111111111111;
		12'b100111010011: color_data = 12'b111111111111;
		12'b100111010100: color_data = 12'b111111111111;
		12'b100111010101: color_data = 12'b111111111111;
		12'b100111010110: color_data = 12'b111111111111;
		12'b100111010111: color_data = 12'b111111111111;
		12'b100111011000: color_data = 12'b111111111111;
		12'b100111011001: color_data = 12'b111111111111;
		12'b100111011010: color_data = 12'b000000000000;
		12'b100111011011: color_data = 12'b111111111111;
		12'b100111011100: color_data = 12'b111111111111;
		12'b100111011101: color_data = 12'b111111111111;
		12'b100111011110: color_data = 12'b111111111111;
		12'b100111011111: color_data = 12'b111111111111;

		12'b100111100000: color_data = 12'b111111111111;
		12'b100111100001: color_data = 12'b111111111111;
		12'b100111100010: color_data = 12'b111111111111;
		12'b100111100011: color_data = 12'b111111111111;
		12'b100111100100: color_data = 12'b000000000000;
		12'b100111100101: color_data = 12'b000000000000;
		12'b100111100110: color_data = 12'b000000000000;
		12'b100111100111: color_data = 12'b000000000000;
		12'b100111101000: color_data = 12'b000000000000;
		12'b100111101001: color_data = 12'b000000000000;
		12'b100111101010: color_data = 12'b000000000000;
		12'b100111101011: color_data = 12'b111111111111;
		12'b100111101100: color_data = 12'b111111111111;
		12'b100111101101: color_data = 12'b111111111111;
		12'b100111101110: color_data = 12'b111111111111;
		12'b100111101111: color_data = 12'b111111111111;

		12'b100111110000: color_data = 12'b111111111111;
		12'b100111110001: color_data = 12'b111111111111;
		12'b100111110010: color_data = 12'b111111111111;
		12'b100111110011: color_data = 12'b111111111111;
		12'b100111110100: color_data = 12'b111111111111;
		12'b100111110101: color_data = 12'b111111111111;
		12'b100111110110: color_data = 12'b111111111111;
		12'b100111110111: color_data = 12'b111111111111;
		12'b100111111000: color_data = 12'b111111111111;
		12'b100111111001: color_data = 12'b111111111111;
		12'b100111111010: color_data = 12'b111111111111;
		12'b100111111011: color_data = 12'b111111111111;
		12'b100111111100: color_data = 12'b111111111111;
		12'b100111111101: color_data = 12'b111111111111;
		12'b100111111110: color_data = 12'b111111111111;
		12'b100111111111: color_data = 12'b111111111111;

		default: color_data = 12'b000000000000;
	endcase
endmodule